magic
tech sky130A
magscale 1 2
timestamp 1709879588
<< checkpaint >>
rect -3418 -3436 35740 26236
<< viali >>
rect 857 21641 891 21675
rect 1593 21641 1627 21675
rect 2329 21641 2363 21675
rect 3249 21641 3283 21675
rect 3801 21641 3835 21675
rect 4537 21641 4571 21675
rect 5273 21641 5307 21675
rect 6009 21641 6043 21675
rect 6745 21641 6779 21675
rect 7481 21641 7515 21675
rect 8401 21641 8435 21675
rect 8953 21641 8987 21675
rect 9689 21641 9723 21675
rect 10425 21641 10459 21675
rect 11161 21641 11195 21675
rect 11897 21641 11931 21675
rect 12633 21641 12667 21675
rect 13553 21641 13587 21675
rect 14105 21641 14139 21675
rect 14841 21641 14875 21675
rect 15577 21641 15611 21675
rect 16313 21641 16347 21675
rect 17049 21641 17083 21675
rect 29009 21641 29043 21675
rect 29561 21641 29595 21675
rect 27169 21505 27203 21539
rect 26985 21437 27019 21471
rect 29193 21437 29227 21471
rect 29745 21437 29779 21471
rect 25973 21369 26007 21403
rect 26801 21369 26835 21403
rect 25697 21301 25731 21335
<< metal1 >>
rect 27154 21904 27160 21956
rect 27212 21944 27218 21956
rect 28994 21944 29000 21956
rect 27212 21916 29000 21944
rect 27212 21904 27218 21916
rect 28994 21904 29000 21916
rect 29052 21904 29058 21956
rect 26970 21836 26976 21888
rect 27028 21876 27034 21888
rect 29546 21876 29552 21888
rect 27028 21848 29552 21876
rect 27028 21836 27034 21848
rect 29546 21836 29552 21848
rect 29604 21836 29610 21888
rect 552 21786 31648 21808
rect 552 21734 4285 21786
rect 4337 21734 4349 21786
rect 4401 21734 4413 21786
rect 4465 21734 4477 21786
rect 4529 21734 4541 21786
rect 4593 21734 12059 21786
rect 12111 21734 12123 21786
rect 12175 21734 12187 21786
rect 12239 21734 12251 21786
rect 12303 21734 12315 21786
rect 12367 21734 19833 21786
rect 19885 21734 19897 21786
rect 19949 21734 19961 21786
rect 20013 21734 20025 21786
rect 20077 21734 20089 21786
rect 20141 21734 27607 21786
rect 27659 21734 27671 21786
rect 27723 21734 27735 21786
rect 27787 21734 27799 21786
rect 27851 21734 27863 21786
rect 27915 21734 31648 21786
rect 552 21712 31648 21734
rect 842 21632 848 21684
rect 900 21632 906 21684
rect 1578 21632 1584 21684
rect 1636 21632 1642 21684
rect 2314 21632 2320 21684
rect 2372 21632 2378 21684
rect 3234 21632 3240 21684
rect 3292 21632 3298 21684
rect 3786 21632 3792 21684
rect 3844 21632 3850 21684
rect 4525 21675 4583 21681
rect 4525 21641 4537 21675
rect 4571 21672 4583 21675
rect 4614 21672 4620 21684
rect 4571 21644 4620 21672
rect 4571 21641 4583 21644
rect 4525 21635 4583 21641
rect 4614 21632 4620 21644
rect 4672 21632 4678 21684
rect 5258 21632 5264 21684
rect 5316 21632 5322 21684
rect 5994 21632 6000 21684
rect 6052 21632 6058 21684
rect 6730 21632 6736 21684
rect 6788 21632 6794 21684
rect 7466 21632 7472 21684
rect 7524 21632 7530 21684
rect 8386 21632 8392 21684
rect 8444 21632 8450 21684
rect 8938 21632 8944 21684
rect 8996 21632 9002 21684
rect 9674 21632 9680 21684
rect 9732 21632 9738 21684
rect 10410 21632 10416 21684
rect 10468 21632 10474 21684
rect 11146 21632 11152 21684
rect 11204 21632 11210 21684
rect 11882 21632 11888 21684
rect 11940 21632 11946 21684
rect 12618 21632 12624 21684
rect 12676 21632 12682 21684
rect 13538 21632 13544 21684
rect 13596 21632 13602 21684
rect 14090 21632 14096 21684
rect 14148 21632 14154 21684
rect 14826 21632 14832 21684
rect 14884 21632 14890 21684
rect 15562 21632 15568 21684
rect 15620 21632 15626 21684
rect 16298 21632 16304 21684
rect 16356 21632 16362 21684
rect 17034 21632 17040 21684
rect 17092 21632 17098 21684
rect 28994 21632 29000 21684
rect 29052 21632 29058 21684
rect 29546 21632 29552 21684
rect 29604 21632 29610 21684
rect 27154 21496 27160 21548
rect 27212 21496 27218 21548
rect 26970 21428 26976 21480
rect 27028 21428 27034 21480
rect 29178 21428 29184 21480
rect 29236 21428 29242 21480
rect 29730 21428 29736 21480
rect 29788 21428 29794 21480
rect 25961 21403 26019 21409
rect 25961 21369 25973 21403
rect 26007 21400 26019 21403
rect 26789 21403 26847 21409
rect 26789 21400 26801 21403
rect 26007 21372 26801 21400
rect 26007 21369 26019 21372
rect 25961 21363 26019 21369
rect 26789 21369 26801 21372
rect 26835 21369 26847 21403
rect 26789 21363 26847 21369
rect 25682 21292 25688 21344
rect 25740 21292 25746 21344
rect 552 21242 31808 21264
rect 552 21190 8172 21242
rect 8224 21190 8236 21242
rect 8288 21190 8300 21242
rect 8352 21190 8364 21242
rect 8416 21190 8428 21242
rect 8480 21190 15946 21242
rect 15998 21190 16010 21242
rect 16062 21190 16074 21242
rect 16126 21190 16138 21242
rect 16190 21190 16202 21242
rect 16254 21190 23720 21242
rect 23772 21190 23784 21242
rect 23836 21190 23848 21242
rect 23900 21190 23912 21242
rect 23964 21190 23976 21242
rect 24028 21190 31494 21242
rect 31546 21190 31558 21242
rect 31610 21190 31622 21242
rect 31674 21190 31686 21242
rect 31738 21190 31750 21242
rect 31802 21190 31808 21242
rect 552 21168 31808 21190
rect 552 20698 31648 20720
rect 552 20646 4285 20698
rect 4337 20646 4349 20698
rect 4401 20646 4413 20698
rect 4465 20646 4477 20698
rect 4529 20646 4541 20698
rect 4593 20646 12059 20698
rect 12111 20646 12123 20698
rect 12175 20646 12187 20698
rect 12239 20646 12251 20698
rect 12303 20646 12315 20698
rect 12367 20646 19833 20698
rect 19885 20646 19897 20698
rect 19949 20646 19961 20698
rect 20013 20646 20025 20698
rect 20077 20646 20089 20698
rect 20141 20646 27607 20698
rect 27659 20646 27671 20698
rect 27723 20646 27735 20698
rect 27787 20646 27799 20698
rect 27851 20646 27863 20698
rect 27915 20646 31648 20698
rect 552 20624 31648 20646
rect 552 20154 31808 20176
rect 552 20102 8172 20154
rect 8224 20102 8236 20154
rect 8288 20102 8300 20154
rect 8352 20102 8364 20154
rect 8416 20102 8428 20154
rect 8480 20102 15946 20154
rect 15998 20102 16010 20154
rect 16062 20102 16074 20154
rect 16126 20102 16138 20154
rect 16190 20102 16202 20154
rect 16254 20102 23720 20154
rect 23772 20102 23784 20154
rect 23836 20102 23848 20154
rect 23900 20102 23912 20154
rect 23964 20102 23976 20154
rect 24028 20102 31494 20154
rect 31546 20102 31558 20154
rect 31610 20102 31622 20154
rect 31674 20102 31686 20154
rect 31738 20102 31750 20154
rect 31802 20102 31808 20154
rect 552 20080 31808 20102
rect 552 19610 31648 19632
rect 552 19558 4285 19610
rect 4337 19558 4349 19610
rect 4401 19558 4413 19610
rect 4465 19558 4477 19610
rect 4529 19558 4541 19610
rect 4593 19558 12059 19610
rect 12111 19558 12123 19610
rect 12175 19558 12187 19610
rect 12239 19558 12251 19610
rect 12303 19558 12315 19610
rect 12367 19558 19833 19610
rect 19885 19558 19897 19610
rect 19949 19558 19961 19610
rect 20013 19558 20025 19610
rect 20077 19558 20089 19610
rect 20141 19558 27607 19610
rect 27659 19558 27671 19610
rect 27723 19558 27735 19610
rect 27787 19558 27799 19610
rect 27851 19558 27863 19610
rect 27915 19558 31648 19610
rect 552 19536 31648 19558
rect 552 19066 31808 19088
rect 552 19014 8172 19066
rect 8224 19014 8236 19066
rect 8288 19014 8300 19066
rect 8352 19014 8364 19066
rect 8416 19014 8428 19066
rect 8480 19014 15946 19066
rect 15998 19014 16010 19066
rect 16062 19014 16074 19066
rect 16126 19014 16138 19066
rect 16190 19014 16202 19066
rect 16254 19014 23720 19066
rect 23772 19014 23784 19066
rect 23836 19014 23848 19066
rect 23900 19014 23912 19066
rect 23964 19014 23976 19066
rect 24028 19014 31494 19066
rect 31546 19014 31558 19066
rect 31610 19014 31622 19066
rect 31674 19014 31686 19066
rect 31738 19014 31750 19066
rect 31802 19014 31808 19066
rect 552 18992 31808 19014
rect 552 18522 31648 18544
rect 552 18470 4285 18522
rect 4337 18470 4349 18522
rect 4401 18470 4413 18522
rect 4465 18470 4477 18522
rect 4529 18470 4541 18522
rect 4593 18470 12059 18522
rect 12111 18470 12123 18522
rect 12175 18470 12187 18522
rect 12239 18470 12251 18522
rect 12303 18470 12315 18522
rect 12367 18470 19833 18522
rect 19885 18470 19897 18522
rect 19949 18470 19961 18522
rect 20013 18470 20025 18522
rect 20077 18470 20089 18522
rect 20141 18470 27607 18522
rect 27659 18470 27671 18522
rect 27723 18470 27735 18522
rect 27787 18470 27799 18522
rect 27851 18470 27863 18522
rect 27915 18470 31648 18522
rect 552 18448 31648 18470
rect 552 17978 31808 18000
rect 552 17926 8172 17978
rect 8224 17926 8236 17978
rect 8288 17926 8300 17978
rect 8352 17926 8364 17978
rect 8416 17926 8428 17978
rect 8480 17926 15946 17978
rect 15998 17926 16010 17978
rect 16062 17926 16074 17978
rect 16126 17926 16138 17978
rect 16190 17926 16202 17978
rect 16254 17926 23720 17978
rect 23772 17926 23784 17978
rect 23836 17926 23848 17978
rect 23900 17926 23912 17978
rect 23964 17926 23976 17978
rect 24028 17926 31494 17978
rect 31546 17926 31558 17978
rect 31610 17926 31622 17978
rect 31674 17926 31686 17978
rect 31738 17926 31750 17978
rect 31802 17926 31808 17978
rect 552 17904 31808 17926
rect 552 17434 31648 17456
rect 552 17382 4285 17434
rect 4337 17382 4349 17434
rect 4401 17382 4413 17434
rect 4465 17382 4477 17434
rect 4529 17382 4541 17434
rect 4593 17382 12059 17434
rect 12111 17382 12123 17434
rect 12175 17382 12187 17434
rect 12239 17382 12251 17434
rect 12303 17382 12315 17434
rect 12367 17382 19833 17434
rect 19885 17382 19897 17434
rect 19949 17382 19961 17434
rect 20013 17382 20025 17434
rect 20077 17382 20089 17434
rect 20141 17382 27607 17434
rect 27659 17382 27671 17434
rect 27723 17382 27735 17434
rect 27787 17382 27799 17434
rect 27851 17382 27863 17434
rect 27915 17382 31648 17434
rect 552 17360 31648 17382
rect 552 16890 31808 16912
rect 552 16838 8172 16890
rect 8224 16838 8236 16890
rect 8288 16838 8300 16890
rect 8352 16838 8364 16890
rect 8416 16838 8428 16890
rect 8480 16838 15946 16890
rect 15998 16838 16010 16890
rect 16062 16838 16074 16890
rect 16126 16838 16138 16890
rect 16190 16838 16202 16890
rect 16254 16838 23720 16890
rect 23772 16838 23784 16890
rect 23836 16838 23848 16890
rect 23900 16838 23912 16890
rect 23964 16838 23976 16890
rect 24028 16838 31494 16890
rect 31546 16838 31558 16890
rect 31610 16838 31622 16890
rect 31674 16838 31686 16890
rect 31738 16838 31750 16890
rect 31802 16838 31808 16890
rect 552 16816 31808 16838
rect 552 16346 31648 16368
rect 552 16294 4285 16346
rect 4337 16294 4349 16346
rect 4401 16294 4413 16346
rect 4465 16294 4477 16346
rect 4529 16294 4541 16346
rect 4593 16294 12059 16346
rect 12111 16294 12123 16346
rect 12175 16294 12187 16346
rect 12239 16294 12251 16346
rect 12303 16294 12315 16346
rect 12367 16294 19833 16346
rect 19885 16294 19897 16346
rect 19949 16294 19961 16346
rect 20013 16294 20025 16346
rect 20077 16294 20089 16346
rect 20141 16294 27607 16346
rect 27659 16294 27671 16346
rect 27723 16294 27735 16346
rect 27787 16294 27799 16346
rect 27851 16294 27863 16346
rect 27915 16294 31648 16346
rect 552 16272 31648 16294
rect 552 15802 31808 15824
rect 552 15750 8172 15802
rect 8224 15750 8236 15802
rect 8288 15750 8300 15802
rect 8352 15750 8364 15802
rect 8416 15750 8428 15802
rect 8480 15750 15946 15802
rect 15998 15750 16010 15802
rect 16062 15750 16074 15802
rect 16126 15750 16138 15802
rect 16190 15750 16202 15802
rect 16254 15750 23720 15802
rect 23772 15750 23784 15802
rect 23836 15750 23848 15802
rect 23900 15750 23912 15802
rect 23964 15750 23976 15802
rect 24028 15750 31494 15802
rect 31546 15750 31558 15802
rect 31610 15750 31622 15802
rect 31674 15750 31686 15802
rect 31738 15750 31750 15802
rect 31802 15750 31808 15802
rect 552 15728 31808 15750
rect 552 15258 31648 15280
rect 552 15206 4285 15258
rect 4337 15206 4349 15258
rect 4401 15206 4413 15258
rect 4465 15206 4477 15258
rect 4529 15206 4541 15258
rect 4593 15206 12059 15258
rect 12111 15206 12123 15258
rect 12175 15206 12187 15258
rect 12239 15206 12251 15258
rect 12303 15206 12315 15258
rect 12367 15206 19833 15258
rect 19885 15206 19897 15258
rect 19949 15206 19961 15258
rect 20013 15206 20025 15258
rect 20077 15206 20089 15258
rect 20141 15206 27607 15258
rect 27659 15206 27671 15258
rect 27723 15206 27735 15258
rect 27787 15206 27799 15258
rect 27851 15206 27863 15258
rect 27915 15206 31648 15258
rect 552 15184 31648 15206
rect 552 14714 31808 14736
rect 552 14662 8172 14714
rect 8224 14662 8236 14714
rect 8288 14662 8300 14714
rect 8352 14662 8364 14714
rect 8416 14662 8428 14714
rect 8480 14662 15946 14714
rect 15998 14662 16010 14714
rect 16062 14662 16074 14714
rect 16126 14662 16138 14714
rect 16190 14662 16202 14714
rect 16254 14662 23720 14714
rect 23772 14662 23784 14714
rect 23836 14662 23848 14714
rect 23900 14662 23912 14714
rect 23964 14662 23976 14714
rect 24028 14662 31494 14714
rect 31546 14662 31558 14714
rect 31610 14662 31622 14714
rect 31674 14662 31686 14714
rect 31738 14662 31750 14714
rect 31802 14662 31808 14714
rect 552 14640 31808 14662
rect 552 14170 31648 14192
rect 552 14118 4285 14170
rect 4337 14118 4349 14170
rect 4401 14118 4413 14170
rect 4465 14118 4477 14170
rect 4529 14118 4541 14170
rect 4593 14118 12059 14170
rect 12111 14118 12123 14170
rect 12175 14118 12187 14170
rect 12239 14118 12251 14170
rect 12303 14118 12315 14170
rect 12367 14118 19833 14170
rect 19885 14118 19897 14170
rect 19949 14118 19961 14170
rect 20013 14118 20025 14170
rect 20077 14118 20089 14170
rect 20141 14118 27607 14170
rect 27659 14118 27671 14170
rect 27723 14118 27735 14170
rect 27787 14118 27799 14170
rect 27851 14118 27863 14170
rect 27915 14118 31648 14170
rect 552 14096 31648 14118
rect 552 13626 31808 13648
rect 552 13574 8172 13626
rect 8224 13574 8236 13626
rect 8288 13574 8300 13626
rect 8352 13574 8364 13626
rect 8416 13574 8428 13626
rect 8480 13574 15946 13626
rect 15998 13574 16010 13626
rect 16062 13574 16074 13626
rect 16126 13574 16138 13626
rect 16190 13574 16202 13626
rect 16254 13574 23720 13626
rect 23772 13574 23784 13626
rect 23836 13574 23848 13626
rect 23900 13574 23912 13626
rect 23964 13574 23976 13626
rect 24028 13574 31494 13626
rect 31546 13574 31558 13626
rect 31610 13574 31622 13626
rect 31674 13574 31686 13626
rect 31738 13574 31750 13626
rect 31802 13574 31808 13626
rect 552 13552 31808 13574
rect 552 13082 31648 13104
rect 552 13030 4285 13082
rect 4337 13030 4349 13082
rect 4401 13030 4413 13082
rect 4465 13030 4477 13082
rect 4529 13030 4541 13082
rect 4593 13030 12059 13082
rect 12111 13030 12123 13082
rect 12175 13030 12187 13082
rect 12239 13030 12251 13082
rect 12303 13030 12315 13082
rect 12367 13030 19833 13082
rect 19885 13030 19897 13082
rect 19949 13030 19961 13082
rect 20013 13030 20025 13082
rect 20077 13030 20089 13082
rect 20141 13030 27607 13082
rect 27659 13030 27671 13082
rect 27723 13030 27735 13082
rect 27787 13030 27799 13082
rect 27851 13030 27863 13082
rect 27915 13030 31648 13082
rect 552 13008 31648 13030
rect 552 12538 31808 12560
rect 552 12486 8172 12538
rect 8224 12486 8236 12538
rect 8288 12486 8300 12538
rect 8352 12486 8364 12538
rect 8416 12486 8428 12538
rect 8480 12486 15946 12538
rect 15998 12486 16010 12538
rect 16062 12486 16074 12538
rect 16126 12486 16138 12538
rect 16190 12486 16202 12538
rect 16254 12486 23720 12538
rect 23772 12486 23784 12538
rect 23836 12486 23848 12538
rect 23900 12486 23912 12538
rect 23964 12486 23976 12538
rect 24028 12486 31494 12538
rect 31546 12486 31558 12538
rect 31610 12486 31622 12538
rect 31674 12486 31686 12538
rect 31738 12486 31750 12538
rect 31802 12486 31808 12538
rect 552 12464 31808 12486
rect 552 11994 31648 12016
rect 552 11942 4285 11994
rect 4337 11942 4349 11994
rect 4401 11942 4413 11994
rect 4465 11942 4477 11994
rect 4529 11942 4541 11994
rect 4593 11942 12059 11994
rect 12111 11942 12123 11994
rect 12175 11942 12187 11994
rect 12239 11942 12251 11994
rect 12303 11942 12315 11994
rect 12367 11942 19833 11994
rect 19885 11942 19897 11994
rect 19949 11942 19961 11994
rect 20013 11942 20025 11994
rect 20077 11942 20089 11994
rect 20141 11942 27607 11994
rect 27659 11942 27671 11994
rect 27723 11942 27735 11994
rect 27787 11942 27799 11994
rect 27851 11942 27863 11994
rect 27915 11942 31648 11994
rect 552 11920 31648 11942
rect 552 11450 31808 11472
rect 552 11398 8172 11450
rect 8224 11398 8236 11450
rect 8288 11398 8300 11450
rect 8352 11398 8364 11450
rect 8416 11398 8428 11450
rect 8480 11398 15946 11450
rect 15998 11398 16010 11450
rect 16062 11398 16074 11450
rect 16126 11398 16138 11450
rect 16190 11398 16202 11450
rect 16254 11398 23720 11450
rect 23772 11398 23784 11450
rect 23836 11398 23848 11450
rect 23900 11398 23912 11450
rect 23964 11398 23976 11450
rect 24028 11398 31494 11450
rect 31546 11398 31558 11450
rect 31610 11398 31622 11450
rect 31674 11398 31686 11450
rect 31738 11398 31750 11450
rect 31802 11398 31808 11450
rect 552 11376 31808 11398
rect 552 10906 31648 10928
rect 552 10854 4285 10906
rect 4337 10854 4349 10906
rect 4401 10854 4413 10906
rect 4465 10854 4477 10906
rect 4529 10854 4541 10906
rect 4593 10854 12059 10906
rect 12111 10854 12123 10906
rect 12175 10854 12187 10906
rect 12239 10854 12251 10906
rect 12303 10854 12315 10906
rect 12367 10854 19833 10906
rect 19885 10854 19897 10906
rect 19949 10854 19961 10906
rect 20013 10854 20025 10906
rect 20077 10854 20089 10906
rect 20141 10854 27607 10906
rect 27659 10854 27671 10906
rect 27723 10854 27735 10906
rect 27787 10854 27799 10906
rect 27851 10854 27863 10906
rect 27915 10854 31648 10906
rect 552 10832 31648 10854
rect 552 10362 31808 10384
rect 552 10310 8172 10362
rect 8224 10310 8236 10362
rect 8288 10310 8300 10362
rect 8352 10310 8364 10362
rect 8416 10310 8428 10362
rect 8480 10310 15946 10362
rect 15998 10310 16010 10362
rect 16062 10310 16074 10362
rect 16126 10310 16138 10362
rect 16190 10310 16202 10362
rect 16254 10310 23720 10362
rect 23772 10310 23784 10362
rect 23836 10310 23848 10362
rect 23900 10310 23912 10362
rect 23964 10310 23976 10362
rect 24028 10310 31494 10362
rect 31546 10310 31558 10362
rect 31610 10310 31622 10362
rect 31674 10310 31686 10362
rect 31738 10310 31750 10362
rect 31802 10310 31808 10362
rect 552 10288 31808 10310
rect 552 9818 31648 9840
rect 552 9766 4285 9818
rect 4337 9766 4349 9818
rect 4401 9766 4413 9818
rect 4465 9766 4477 9818
rect 4529 9766 4541 9818
rect 4593 9766 12059 9818
rect 12111 9766 12123 9818
rect 12175 9766 12187 9818
rect 12239 9766 12251 9818
rect 12303 9766 12315 9818
rect 12367 9766 19833 9818
rect 19885 9766 19897 9818
rect 19949 9766 19961 9818
rect 20013 9766 20025 9818
rect 20077 9766 20089 9818
rect 20141 9766 27607 9818
rect 27659 9766 27671 9818
rect 27723 9766 27735 9818
rect 27787 9766 27799 9818
rect 27851 9766 27863 9818
rect 27915 9766 31648 9818
rect 552 9744 31648 9766
rect 552 9274 31808 9296
rect 552 9222 8172 9274
rect 8224 9222 8236 9274
rect 8288 9222 8300 9274
rect 8352 9222 8364 9274
rect 8416 9222 8428 9274
rect 8480 9222 15946 9274
rect 15998 9222 16010 9274
rect 16062 9222 16074 9274
rect 16126 9222 16138 9274
rect 16190 9222 16202 9274
rect 16254 9222 23720 9274
rect 23772 9222 23784 9274
rect 23836 9222 23848 9274
rect 23900 9222 23912 9274
rect 23964 9222 23976 9274
rect 24028 9222 31494 9274
rect 31546 9222 31558 9274
rect 31610 9222 31622 9274
rect 31674 9222 31686 9274
rect 31738 9222 31750 9274
rect 31802 9222 31808 9274
rect 552 9200 31808 9222
rect 552 8730 31648 8752
rect 552 8678 4285 8730
rect 4337 8678 4349 8730
rect 4401 8678 4413 8730
rect 4465 8678 4477 8730
rect 4529 8678 4541 8730
rect 4593 8678 12059 8730
rect 12111 8678 12123 8730
rect 12175 8678 12187 8730
rect 12239 8678 12251 8730
rect 12303 8678 12315 8730
rect 12367 8678 19833 8730
rect 19885 8678 19897 8730
rect 19949 8678 19961 8730
rect 20013 8678 20025 8730
rect 20077 8678 20089 8730
rect 20141 8678 27607 8730
rect 27659 8678 27671 8730
rect 27723 8678 27735 8730
rect 27787 8678 27799 8730
rect 27851 8678 27863 8730
rect 27915 8678 31648 8730
rect 552 8656 31648 8678
rect 552 8186 31808 8208
rect 552 8134 8172 8186
rect 8224 8134 8236 8186
rect 8288 8134 8300 8186
rect 8352 8134 8364 8186
rect 8416 8134 8428 8186
rect 8480 8134 15946 8186
rect 15998 8134 16010 8186
rect 16062 8134 16074 8186
rect 16126 8134 16138 8186
rect 16190 8134 16202 8186
rect 16254 8134 23720 8186
rect 23772 8134 23784 8186
rect 23836 8134 23848 8186
rect 23900 8134 23912 8186
rect 23964 8134 23976 8186
rect 24028 8134 31494 8186
rect 31546 8134 31558 8186
rect 31610 8134 31622 8186
rect 31674 8134 31686 8186
rect 31738 8134 31750 8186
rect 31802 8134 31808 8186
rect 552 8112 31808 8134
rect 552 7642 31648 7664
rect 552 7590 4285 7642
rect 4337 7590 4349 7642
rect 4401 7590 4413 7642
rect 4465 7590 4477 7642
rect 4529 7590 4541 7642
rect 4593 7590 12059 7642
rect 12111 7590 12123 7642
rect 12175 7590 12187 7642
rect 12239 7590 12251 7642
rect 12303 7590 12315 7642
rect 12367 7590 19833 7642
rect 19885 7590 19897 7642
rect 19949 7590 19961 7642
rect 20013 7590 20025 7642
rect 20077 7590 20089 7642
rect 20141 7590 27607 7642
rect 27659 7590 27671 7642
rect 27723 7590 27735 7642
rect 27787 7590 27799 7642
rect 27851 7590 27863 7642
rect 27915 7590 31648 7642
rect 552 7568 31648 7590
rect 552 7098 31808 7120
rect 552 7046 8172 7098
rect 8224 7046 8236 7098
rect 8288 7046 8300 7098
rect 8352 7046 8364 7098
rect 8416 7046 8428 7098
rect 8480 7046 15946 7098
rect 15998 7046 16010 7098
rect 16062 7046 16074 7098
rect 16126 7046 16138 7098
rect 16190 7046 16202 7098
rect 16254 7046 23720 7098
rect 23772 7046 23784 7098
rect 23836 7046 23848 7098
rect 23900 7046 23912 7098
rect 23964 7046 23976 7098
rect 24028 7046 31494 7098
rect 31546 7046 31558 7098
rect 31610 7046 31622 7098
rect 31674 7046 31686 7098
rect 31738 7046 31750 7098
rect 31802 7046 31808 7098
rect 552 7024 31808 7046
rect 552 6554 31648 6576
rect 552 6502 4285 6554
rect 4337 6502 4349 6554
rect 4401 6502 4413 6554
rect 4465 6502 4477 6554
rect 4529 6502 4541 6554
rect 4593 6502 12059 6554
rect 12111 6502 12123 6554
rect 12175 6502 12187 6554
rect 12239 6502 12251 6554
rect 12303 6502 12315 6554
rect 12367 6502 19833 6554
rect 19885 6502 19897 6554
rect 19949 6502 19961 6554
rect 20013 6502 20025 6554
rect 20077 6502 20089 6554
rect 20141 6502 27607 6554
rect 27659 6502 27671 6554
rect 27723 6502 27735 6554
rect 27787 6502 27799 6554
rect 27851 6502 27863 6554
rect 27915 6502 31648 6554
rect 552 6480 31648 6502
rect 552 6010 31808 6032
rect 552 5958 8172 6010
rect 8224 5958 8236 6010
rect 8288 5958 8300 6010
rect 8352 5958 8364 6010
rect 8416 5958 8428 6010
rect 8480 5958 15946 6010
rect 15998 5958 16010 6010
rect 16062 5958 16074 6010
rect 16126 5958 16138 6010
rect 16190 5958 16202 6010
rect 16254 5958 23720 6010
rect 23772 5958 23784 6010
rect 23836 5958 23848 6010
rect 23900 5958 23912 6010
rect 23964 5958 23976 6010
rect 24028 5958 31494 6010
rect 31546 5958 31558 6010
rect 31610 5958 31622 6010
rect 31674 5958 31686 6010
rect 31738 5958 31750 6010
rect 31802 5958 31808 6010
rect 552 5936 31808 5958
rect 552 5466 31648 5488
rect 552 5414 4285 5466
rect 4337 5414 4349 5466
rect 4401 5414 4413 5466
rect 4465 5414 4477 5466
rect 4529 5414 4541 5466
rect 4593 5414 12059 5466
rect 12111 5414 12123 5466
rect 12175 5414 12187 5466
rect 12239 5414 12251 5466
rect 12303 5414 12315 5466
rect 12367 5414 19833 5466
rect 19885 5414 19897 5466
rect 19949 5414 19961 5466
rect 20013 5414 20025 5466
rect 20077 5414 20089 5466
rect 20141 5414 27607 5466
rect 27659 5414 27671 5466
rect 27723 5414 27735 5466
rect 27787 5414 27799 5466
rect 27851 5414 27863 5466
rect 27915 5414 31648 5466
rect 552 5392 31648 5414
rect 552 4922 31808 4944
rect 552 4870 8172 4922
rect 8224 4870 8236 4922
rect 8288 4870 8300 4922
rect 8352 4870 8364 4922
rect 8416 4870 8428 4922
rect 8480 4870 15946 4922
rect 15998 4870 16010 4922
rect 16062 4870 16074 4922
rect 16126 4870 16138 4922
rect 16190 4870 16202 4922
rect 16254 4870 23720 4922
rect 23772 4870 23784 4922
rect 23836 4870 23848 4922
rect 23900 4870 23912 4922
rect 23964 4870 23976 4922
rect 24028 4870 31494 4922
rect 31546 4870 31558 4922
rect 31610 4870 31622 4922
rect 31674 4870 31686 4922
rect 31738 4870 31750 4922
rect 31802 4870 31808 4922
rect 552 4848 31808 4870
rect 552 4378 31648 4400
rect 552 4326 4285 4378
rect 4337 4326 4349 4378
rect 4401 4326 4413 4378
rect 4465 4326 4477 4378
rect 4529 4326 4541 4378
rect 4593 4326 12059 4378
rect 12111 4326 12123 4378
rect 12175 4326 12187 4378
rect 12239 4326 12251 4378
rect 12303 4326 12315 4378
rect 12367 4326 19833 4378
rect 19885 4326 19897 4378
rect 19949 4326 19961 4378
rect 20013 4326 20025 4378
rect 20077 4326 20089 4378
rect 20141 4326 27607 4378
rect 27659 4326 27671 4378
rect 27723 4326 27735 4378
rect 27787 4326 27799 4378
rect 27851 4326 27863 4378
rect 27915 4326 31648 4378
rect 552 4304 31648 4326
rect 552 3834 31808 3856
rect 552 3782 8172 3834
rect 8224 3782 8236 3834
rect 8288 3782 8300 3834
rect 8352 3782 8364 3834
rect 8416 3782 8428 3834
rect 8480 3782 15946 3834
rect 15998 3782 16010 3834
rect 16062 3782 16074 3834
rect 16126 3782 16138 3834
rect 16190 3782 16202 3834
rect 16254 3782 23720 3834
rect 23772 3782 23784 3834
rect 23836 3782 23848 3834
rect 23900 3782 23912 3834
rect 23964 3782 23976 3834
rect 24028 3782 31494 3834
rect 31546 3782 31558 3834
rect 31610 3782 31622 3834
rect 31674 3782 31686 3834
rect 31738 3782 31750 3834
rect 31802 3782 31808 3834
rect 552 3760 31808 3782
rect 552 3290 31648 3312
rect 552 3238 4285 3290
rect 4337 3238 4349 3290
rect 4401 3238 4413 3290
rect 4465 3238 4477 3290
rect 4529 3238 4541 3290
rect 4593 3238 12059 3290
rect 12111 3238 12123 3290
rect 12175 3238 12187 3290
rect 12239 3238 12251 3290
rect 12303 3238 12315 3290
rect 12367 3238 19833 3290
rect 19885 3238 19897 3290
rect 19949 3238 19961 3290
rect 20013 3238 20025 3290
rect 20077 3238 20089 3290
rect 20141 3238 27607 3290
rect 27659 3238 27671 3290
rect 27723 3238 27735 3290
rect 27787 3238 27799 3290
rect 27851 3238 27863 3290
rect 27915 3238 31648 3290
rect 552 3216 31648 3238
rect 552 2746 31808 2768
rect 552 2694 8172 2746
rect 8224 2694 8236 2746
rect 8288 2694 8300 2746
rect 8352 2694 8364 2746
rect 8416 2694 8428 2746
rect 8480 2694 15946 2746
rect 15998 2694 16010 2746
rect 16062 2694 16074 2746
rect 16126 2694 16138 2746
rect 16190 2694 16202 2746
rect 16254 2694 23720 2746
rect 23772 2694 23784 2746
rect 23836 2694 23848 2746
rect 23900 2694 23912 2746
rect 23964 2694 23976 2746
rect 24028 2694 31494 2746
rect 31546 2694 31558 2746
rect 31610 2694 31622 2746
rect 31674 2694 31686 2746
rect 31738 2694 31750 2746
rect 31802 2694 31808 2746
rect 552 2672 31808 2694
rect 552 2202 31648 2224
rect 552 2150 4285 2202
rect 4337 2150 4349 2202
rect 4401 2150 4413 2202
rect 4465 2150 4477 2202
rect 4529 2150 4541 2202
rect 4593 2150 12059 2202
rect 12111 2150 12123 2202
rect 12175 2150 12187 2202
rect 12239 2150 12251 2202
rect 12303 2150 12315 2202
rect 12367 2150 19833 2202
rect 19885 2150 19897 2202
rect 19949 2150 19961 2202
rect 20013 2150 20025 2202
rect 20077 2150 20089 2202
rect 20141 2150 27607 2202
rect 27659 2150 27671 2202
rect 27723 2150 27735 2202
rect 27787 2150 27799 2202
rect 27851 2150 27863 2202
rect 27915 2150 31648 2202
rect 552 2128 31648 2150
rect 552 1658 31808 1680
rect 552 1606 8172 1658
rect 8224 1606 8236 1658
rect 8288 1606 8300 1658
rect 8352 1606 8364 1658
rect 8416 1606 8428 1658
rect 8480 1606 15946 1658
rect 15998 1606 16010 1658
rect 16062 1606 16074 1658
rect 16126 1606 16138 1658
rect 16190 1606 16202 1658
rect 16254 1606 23720 1658
rect 23772 1606 23784 1658
rect 23836 1606 23848 1658
rect 23900 1606 23912 1658
rect 23964 1606 23976 1658
rect 24028 1606 31494 1658
rect 31546 1606 31558 1658
rect 31610 1606 31622 1658
rect 31674 1606 31686 1658
rect 31738 1606 31750 1658
rect 31802 1606 31808 1658
rect 552 1584 31808 1606
rect 552 1114 31648 1136
rect 552 1062 4285 1114
rect 4337 1062 4349 1114
rect 4401 1062 4413 1114
rect 4465 1062 4477 1114
rect 4529 1062 4541 1114
rect 4593 1062 12059 1114
rect 12111 1062 12123 1114
rect 12175 1062 12187 1114
rect 12239 1062 12251 1114
rect 12303 1062 12315 1114
rect 12367 1062 19833 1114
rect 19885 1062 19897 1114
rect 19949 1062 19961 1114
rect 20013 1062 20025 1114
rect 20077 1062 20089 1114
rect 20141 1062 27607 1114
rect 27659 1062 27671 1114
rect 27723 1062 27735 1114
rect 27787 1062 27799 1114
rect 27851 1062 27863 1114
rect 27915 1062 31648 1114
rect 552 1040 31648 1062
rect 552 570 31808 592
rect 552 518 8172 570
rect 8224 518 8236 570
rect 8288 518 8300 570
rect 8352 518 8364 570
rect 8416 518 8428 570
rect 8480 518 15946 570
rect 15998 518 16010 570
rect 16062 518 16074 570
rect 16126 518 16138 570
rect 16190 518 16202 570
rect 16254 518 23720 570
rect 23772 518 23784 570
rect 23836 518 23848 570
rect 23900 518 23912 570
rect 23964 518 23976 570
rect 24028 518 31494 570
rect 31546 518 31558 570
rect 31610 518 31622 570
rect 31674 518 31686 570
rect 31738 518 31750 570
rect 31802 518 31808 570
rect 552 496 31808 518
<< via1 >>
rect 27160 21904 27212 21956
rect 29000 21904 29052 21956
rect 26976 21836 27028 21888
rect 29552 21836 29604 21888
rect 4285 21734 4337 21786
rect 4349 21734 4401 21786
rect 4413 21734 4465 21786
rect 4477 21734 4529 21786
rect 4541 21734 4593 21786
rect 12059 21734 12111 21786
rect 12123 21734 12175 21786
rect 12187 21734 12239 21786
rect 12251 21734 12303 21786
rect 12315 21734 12367 21786
rect 19833 21734 19885 21786
rect 19897 21734 19949 21786
rect 19961 21734 20013 21786
rect 20025 21734 20077 21786
rect 20089 21734 20141 21786
rect 27607 21734 27659 21786
rect 27671 21734 27723 21786
rect 27735 21734 27787 21786
rect 27799 21734 27851 21786
rect 27863 21734 27915 21786
rect 848 21675 900 21684
rect 848 21641 857 21675
rect 857 21641 891 21675
rect 891 21641 900 21675
rect 848 21632 900 21641
rect 1584 21675 1636 21684
rect 1584 21641 1593 21675
rect 1593 21641 1627 21675
rect 1627 21641 1636 21675
rect 1584 21632 1636 21641
rect 2320 21675 2372 21684
rect 2320 21641 2329 21675
rect 2329 21641 2363 21675
rect 2363 21641 2372 21675
rect 2320 21632 2372 21641
rect 3240 21675 3292 21684
rect 3240 21641 3249 21675
rect 3249 21641 3283 21675
rect 3283 21641 3292 21675
rect 3240 21632 3292 21641
rect 3792 21675 3844 21684
rect 3792 21641 3801 21675
rect 3801 21641 3835 21675
rect 3835 21641 3844 21675
rect 3792 21632 3844 21641
rect 4620 21632 4672 21684
rect 5264 21675 5316 21684
rect 5264 21641 5273 21675
rect 5273 21641 5307 21675
rect 5307 21641 5316 21675
rect 5264 21632 5316 21641
rect 6000 21675 6052 21684
rect 6000 21641 6009 21675
rect 6009 21641 6043 21675
rect 6043 21641 6052 21675
rect 6000 21632 6052 21641
rect 6736 21675 6788 21684
rect 6736 21641 6745 21675
rect 6745 21641 6779 21675
rect 6779 21641 6788 21675
rect 6736 21632 6788 21641
rect 7472 21675 7524 21684
rect 7472 21641 7481 21675
rect 7481 21641 7515 21675
rect 7515 21641 7524 21675
rect 7472 21632 7524 21641
rect 8392 21675 8444 21684
rect 8392 21641 8401 21675
rect 8401 21641 8435 21675
rect 8435 21641 8444 21675
rect 8392 21632 8444 21641
rect 8944 21675 8996 21684
rect 8944 21641 8953 21675
rect 8953 21641 8987 21675
rect 8987 21641 8996 21675
rect 8944 21632 8996 21641
rect 9680 21675 9732 21684
rect 9680 21641 9689 21675
rect 9689 21641 9723 21675
rect 9723 21641 9732 21675
rect 9680 21632 9732 21641
rect 10416 21675 10468 21684
rect 10416 21641 10425 21675
rect 10425 21641 10459 21675
rect 10459 21641 10468 21675
rect 10416 21632 10468 21641
rect 11152 21675 11204 21684
rect 11152 21641 11161 21675
rect 11161 21641 11195 21675
rect 11195 21641 11204 21675
rect 11152 21632 11204 21641
rect 11888 21675 11940 21684
rect 11888 21641 11897 21675
rect 11897 21641 11931 21675
rect 11931 21641 11940 21675
rect 11888 21632 11940 21641
rect 12624 21675 12676 21684
rect 12624 21641 12633 21675
rect 12633 21641 12667 21675
rect 12667 21641 12676 21675
rect 12624 21632 12676 21641
rect 13544 21675 13596 21684
rect 13544 21641 13553 21675
rect 13553 21641 13587 21675
rect 13587 21641 13596 21675
rect 13544 21632 13596 21641
rect 14096 21675 14148 21684
rect 14096 21641 14105 21675
rect 14105 21641 14139 21675
rect 14139 21641 14148 21675
rect 14096 21632 14148 21641
rect 14832 21675 14884 21684
rect 14832 21641 14841 21675
rect 14841 21641 14875 21675
rect 14875 21641 14884 21675
rect 14832 21632 14884 21641
rect 15568 21675 15620 21684
rect 15568 21641 15577 21675
rect 15577 21641 15611 21675
rect 15611 21641 15620 21675
rect 15568 21632 15620 21641
rect 16304 21675 16356 21684
rect 16304 21641 16313 21675
rect 16313 21641 16347 21675
rect 16347 21641 16356 21675
rect 16304 21632 16356 21641
rect 17040 21675 17092 21684
rect 17040 21641 17049 21675
rect 17049 21641 17083 21675
rect 17083 21641 17092 21675
rect 17040 21632 17092 21641
rect 29000 21675 29052 21684
rect 29000 21641 29009 21675
rect 29009 21641 29043 21675
rect 29043 21641 29052 21675
rect 29000 21632 29052 21641
rect 29552 21675 29604 21684
rect 29552 21641 29561 21675
rect 29561 21641 29595 21675
rect 29595 21641 29604 21675
rect 29552 21632 29604 21641
rect 27160 21539 27212 21548
rect 27160 21505 27169 21539
rect 27169 21505 27203 21539
rect 27203 21505 27212 21539
rect 27160 21496 27212 21505
rect 26976 21471 27028 21480
rect 26976 21437 26985 21471
rect 26985 21437 27019 21471
rect 27019 21437 27028 21471
rect 26976 21428 27028 21437
rect 29184 21471 29236 21480
rect 29184 21437 29193 21471
rect 29193 21437 29227 21471
rect 29227 21437 29236 21471
rect 29184 21428 29236 21437
rect 29736 21471 29788 21480
rect 29736 21437 29745 21471
rect 29745 21437 29779 21471
rect 29779 21437 29788 21471
rect 29736 21428 29788 21437
rect 25688 21335 25740 21344
rect 25688 21301 25697 21335
rect 25697 21301 25731 21335
rect 25731 21301 25740 21335
rect 25688 21292 25740 21301
rect 8172 21190 8224 21242
rect 8236 21190 8288 21242
rect 8300 21190 8352 21242
rect 8364 21190 8416 21242
rect 8428 21190 8480 21242
rect 15946 21190 15998 21242
rect 16010 21190 16062 21242
rect 16074 21190 16126 21242
rect 16138 21190 16190 21242
rect 16202 21190 16254 21242
rect 23720 21190 23772 21242
rect 23784 21190 23836 21242
rect 23848 21190 23900 21242
rect 23912 21190 23964 21242
rect 23976 21190 24028 21242
rect 31494 21190 31546 21242
rect 31558 21190 31610 21242
rect 31622 21190 31674 21242
rect 31686 21190 31738 21242
rect 31750 21190 31802 21242
rect 4285 20646 4337 20698
rect 4349 20646 4401 20698
rect 4413 20646 4465 20698
rect 4477 20646 4529 20698
rect 4541 20646 4593 20698
rect 12059 20646 12111 20698
rect 12123 20646 12175 20698
rect 12187 20646 12239 20698
rect 12251 20646 12303 20698
rect 12315 20646 12367 20698
rect 19833 20646 19885 20698
rect 19897 20646 19949 20698
rect 19961 20646 20013 20698
rect 20025 20646 20077 20698
rect 20089 20646 20141 20698
rect 27607 20646 27659 20698
rect 27671 20646 27723 20698
rect 27735 20646 27787 20698
rect 27799 20646 27851 20698
rect 27863 20646 27915 20698
rect 8172 20102 8224 20154
rect 8236 20102 8288 20154
rect 8300 20102 8352 20154
rect 8364 20102 8416 20154
rect 8428 20102 8480 20154
rect 15946 20102 15998 20154
rect 16010 20102 16062 20154
rect 16074 20102 16126 20154
rect 16138 20102 16190 20154
rect 16202 20102 16254 20154
rect 23720 20102 23772 20154
rect 23784 20102 23836 20154
rect 23848 20102 23900 20154
rect 23912 20102 23964 20154
rect 23976 20102 24028 20154
rect 31494 20102 31546 20154
rect 31558 20102 31610 20154
rect 31622 20102 31674 20154
rect 31686 20102 31738 20154
rect 31750 20102 31802 20154
rect 4285 19558 4337 19610
rect 4349 19558 4401 19610
rect 4413 19558 4465 19610
rect 4477 19558 4529 19610
rect 4541 19558 4593 19610
rect 12059 19558 12111 19610
rect 12123 19558 12175 19610
rect 12187 19558 12239 19610
rect 12251 19558 12303 19610
rect 12315 19558 12367 19610
rect 19833 19558 19885 19610
rect 19897 19558 19949 19610
rect 19961 19558 20013 19610
rect 20025 19558 20077 19610
rect 20089 19558 20141 19610
rect 27607 19558 27659 19610
rect 27671 19558 27723 19610
rect 27735 19558 27787 19610
rect 27799 19558 27851 19610
rect 27863 19558 27915 19610
rect 8172 19014 8224 19066
rect 8236 19014 8288 19066
rect 8300 19014 8352 19066
rect 8364 19014 8416 19066
rect 8428 19014 8480 19066
rect 15946 19014 15998 19066
rect 16010 19014 16062 19066
rect 16074 19014 16126 19066
rect 16138 19014 16190 19066
rect 16202 19014 16254 19066
rect 23720 19014 23772 19066
rect 23784 19014 23836 19066
rect 23848 19014 23900 19066
rect 23912 19014 23964 19066
rect 23976 19014 24028 19066
rect 31494 19014 31546 19066
rect 31558 19014 31610 19066
rect 31622 19014 31674 19066
rect 31686 19014 31738 19066
rect 31750 19014 31802 19066
rect 4285 18470 4337 18522
rect 4349 18470 4401 18522
rect 4413 18470 4465 18522
rect 4477 18470 4529 18522
rect 4541 18470 4593 18522
rect 12059 18470 12111 18522
rect 12123 18470 12175 18522
rect 12187 18470 12239 18522
rect 12251 18470 12303 18522
rect 12315 18470 12367 18522
rect 19833 18470 19885 18522
rect 19897 18470 19949 18522
rect 19961 18470 20013 18522
rect 20025 18470 20077 18522
rect 20089 18470 20141 18522
rect 27607 18470 27659 18522
rect 27671 18470 27723 18522
rect 27735 18470 27787 18522
rect 27799 18470 27851 18522
rect 27863 18470 27915 18522
rect 8172 17926 8224 17978
rect 8236 17926 8288 17978
rect 8300 17926 8352 17978
rect 8364 17926 8416 17978
rect 8428 17926 8480 17978
rect 15946 17926 15998 17978
rect 16010 17926 16062 17978
rect 16074 17926 16126 17978
rect 16138 17926 16190 17978
rect 16202 17926 16254 17978
rect 23720 17926 23772 17978
rect 23784 17926 23836 17978
rect 23848 17926 23900 17978
rect 23912 17926 23964 17978
rect 23976 17926 24028 17978
rect 31494 17926 31546 17978
rect 31558 17926 31610 17978
rect 31622 17926 31674 17978
rect 31686 17926 31738 17978
rect 31750 17926 31802 17978
rect 4285 17382 4337 17434
rect 4349 17382 4401 17434
rect 4413 17382 4465 17434
rect 4477 17382 4529 17434
rect 4541 17382 4593 17434
rect 12059 17382 12111 17434
rect 12123 17382 12175 17434
rect 12187 17382 12239 17434
rect 12251 17382 12303 17434
rect 12315 17382 12367 17434
rect 19833 17382 19885 17434
rect 19897 17382 19949 17434
rect 19961 17382 20013 17434
rect 20025 17382 20077 17434
rect 20089 17382 20141 17434
rect 27607 17382 27659 17434
rect 27671 17382 27723 17434
rect 27735 17382 27787 17434
rect 27799 17382 27851 17434
rect 27863 17382 27915 17434
rect 8172 16838 8224 16890
rect 8236 16838 8288 16890
rect 8300 16838 8352 16890
rect 8364 16838 8416 16890
rect 8428 16838 8480 16890
rect 15946 16838 15998 16890
rect 16010 16838 16062 16890
rect 16074 16838 16126 16890
rect 16138 16838 16190 16890
rect 16202 16838 16254 16890
rect 23720 16838 23772 16890
rect 23784 16838 23836 16890
rect 23848 16838 23900 16890
rect 23912 16838 23964 16890
rect 23976 16838 24028 16890
rect 31494 16838 31546 16890
rect 31558 16838 31610 16890
rect 31622 16838 31674 16890
rect 31686 16838 31738 16890
rect 31750 16838 31802 16890
rect 4285 16294 4337 16346
rect 4349 16294 4401 16346
rect 4413 16294 4465 16346
rect 4477 16294 4529 16346
rect 4541 16294 4593 16346
rect 12059 16294 12111 16346
rect 12123 16294 12175 16346
rect 12187 16294 12239 16346
rect 12251 16294 12303 16346
rect 12315 16294 12367 16346
rect 19833 16294 19885 16346
rect 19897 16294 19949 16346
rect 19961 16294 20013 16346
rect 20025 16294 20077 16346
rect 20089 16294 20141 16346
rect 27607 16294 27659 16346
rect 27671 16294 27723 16346
rect 27735 16294 27787 16346
rect 27799 16294 27851 16346
rect 27863 16294 27915 16346
rect 8172 15750 8224 15802
rect 8236 15750 8288 15802
rect 8300 15750 8352 15802
rect 8364 15750 8416 15802
rect 8428 15750 8480 15802
rect 15946 15750 15998 15802
rect 16010 15750 16062 15802
rect 16074 15750 16126 15802
rect 16138 15750 16190 15802
rect 16202 15750 16254 15802
rect 23720 15750 23772 15802
rect 23784 15750 23836 15802
rect 23848 15750 23900 15802
rect 23912 15750 23964 15802
rect 23976 15750 24028 15802
rect 31494 15750 31546 15802
rect 31558 15750 31610 15802
rect 31622 15750 31674 15802
rect 31686 15750 31738 15802
rect 31750 15750 31802 15802
rect 4285 15206 4337 15258
rect 4349 15206 4401 15258
rect 4413 15206 4465 15258
rect 4477 15206 4529 15258
rect 4541 15206 4593 15258
rect 12059 15206 12111 15258
rect 12123 15206 12175 15258
rect 12187 15206 12239 15258
rect 12251 15206 12303 15258
rect 12315 15206 12367 15258
rect 19833 15206 19885 15258
rect 19897 15206 19949 15258
rect 19961 15206 20013 15258
rect 20025 15206 20077 15258
rect 20089 15206 20141 15258
rect 27607 15206 27659 15258
rect 27671 15206 27723 15258
rect 27735 15206 27787 15258
rect 27799 15206 27851 15258
rect 27863 15206 27915 15258
rect 8172 14662 8224 14714
rect 8236 14662 8288 14714
rect 8300 14662 8352 14714
rect 8364 14662 8416 14714
rect 8428 14662 8480 14714
rect 15946 14662 15998 14714
rect 16010 14662 16062 14714
rect 16074 14662 16126 14714
rect 16138 14662 16190 14714
rect 16202 14662 16254 14714
rect 23720 14662 23772 14714
rect 23784 14662 23836 14714
rect 23848 14662 23900 14714
rect 23912 14662 23964 14714
rect 23976 14662 24028 14714
rect 31494 14662 31546 14714
rect 31558 14662 31610 14714
rect 31622 14662 31674 14714
rect 31686 14662 31738 14714
rect 31750 14662 31802 14714
rect 4285 14118 4337 14170
rect 4349 14118 4401 14170
rect 4413 14118 4465 14170
rect 4477 14118 4529 14170
rect 4541 14118 4593 14170
rect 12059 14118 12111 14170
rect 12123 14118 12175 14170
rect 12187 14118 12239 14170
rect 12251 14118 12303 14170
rect 12315 14118 12367 14170
rect 19833 14118 19885 14170
rect 19897 14118 19949 14170
rect 19961 14118 20013 14170
rect 20025 14118 20077 14170
rect 20089 14118 20141 14170
rect 27607 14118 27659 14170
rect 27671 14118 27723 14170
rect 27735 14118 27787 14170
rect 27799 14118 27851 14170
rect 27863 14118 27915 14170
rect 8172 13574 8224 13626
rect 8236 13574 8288 13626
rect 8300 13574 8352 13626
rect 8364 13574 8416 13626
rect 8428 13574 8480 13626
rect 15946 13574 15998 13626
rect 16010 13574 16062 13626
rect 16074 13574 16126 13626
rect 16138 13574 16190 13626
rect 16202 13574 16254 13626
rect 23720 13574 23772 13626
rect 23784 13574 23836 13626
rect 23848 13574 23900 13626
rect 23912 13574 23964 13626
rect 23976 13574 24028 13626
rect 31494 13574 31546 13626
rect 31558 13574 31610 13626
rect 31622 13574 31674 13626
rect 31686 13574 31738 13626
rect 31750 13574 31802 13626
rect 4285 13030 4337 13082
rect 4349 13030 4401 13082
rect 4413 13030 4465 13082
rect 4477 13030 4529 13082
rect 4541 13030 4593 13082
rect 12059 13030 12111 13082
rect 12123 13030 12175 13082
rect 12187 13030 12239 13082
rect 12251 13030 12303 13082
rect 12315 13030 12367 13082
rect 19833 13030 19885 13082
rect 19897 13030 19949 13082
rect 19961 13030 20013 13082
rect 20025 13030 20077 13082
rect 20089 13030 20141 13082
rect 27607 13030 27659 13082
rect 27671 13030 27723 13082
rect 27735 13030 27787 13082
rect 27799 13030 27851 13082
rect 27863 13030 27915 13082
rect 8172 12486 8224 12538
rect 8236 12486 8288 12538
rect 8300 12486 8352 12538
rect 8364 12486 8416 12538
rect 8428 12486 8480 12538
rect 15946 12486 15998 12538
rect 16010 12486 16062 12538
rect 16074 12486 16126 12538
rect 16138 12486 16190 12538
rect 16202 12486 16254 12538
rect 23720 12486 23772 12538
rect 23784 12486 23836 12538
rect 23848 12486 23900 12538
rect 23912 12486 23964 12538
rect 23976 12486 24028 12538
rect 31494 12486 31546 12538
rect 31558 12486 31610 12538
rect 31622 12486 31674 12538
rect 31686 12486 31738 12538
rect 31750 12486 31802 12538
rect 4285 11942 4337 11994
rect 4349 11942 4401 11994
rect 4413 11942 4465 11994
rect 4477 11942 4529 11994
rect 4541 11942 4593 11994
rect 12059 11942 12111 11994
rect 12123 11942 12175 11994
rect 12187 11942 12239 11994
rect 12251 11942 12303 11994
rect 12315 11942 12367 11994
rect 19833 11942 19885 11994
rect 19897 11942 19949 11994
rect 19961 11942 20013 11994
rect 20025 11942 20077 11994
rect 20089 11942 20141 11994
rect 27607 11942 27659 11994
rect 27671 11942 27723 11994
rect 27735 11942 27787 11994
rect 27799 11942 27851 11994
rect 27863 11942 27915 11994
rect 8172 11398 8224 11450
rect 8236 11398 8288 11450
rect 8300 11398 8352 11450
rect 8364 11398 8416 11450
rect 8428 11398 8480 11450
rect 15946 11398 15998 11450
rect 16010 11398 16062 11450
rect 16074 11398 16126 11450
rect 16138 11398 16190 11450
rect 16202 11398 16254 11450
rect 23720 11398 23772 11450
rect 23784 11398 23836 11450
rect 23848 11398 23900 11450
rect 23912 11398 23964 11450
rect 23976 11398 24028 11450
rect 31494 11398 31546 11450
rect 31558 11398 31610 11450
rect 31622 11398 31674 11450
rect 31686 11398 31738 11450
rect 31750 11398 31802 11450
rect 4285 10854 4337 10906
rect 4349 10854 4401 10906
rect 4413 10854 4465 10906
rect 4477 10854 4529 10906
rect 4541 10854 4593 10906
rect 12059 10854 12111 10906
rect 12123 10854 12175 10906
rect 12187 10854 12239 10906
rect 12251 10854 12303 10906
rect 12315 10854 12367 10906
rect 19833 10854 19885 10906
rect 19897 10854 19949 10906
rect 19961 10854 20013 10906
rect 20025 10854 20077 10906
rect 20089 10854 20141 10906
rect 27607 10854 27659 10906
rect 27671 10854 27723 10906
rect 27735 10854 27787 10906
rect 27799 10854 27851 10906
rect 27863 10854 27915 10906
rect 8172 10310 8224 10362
rect 8236 10310 8288 10362
rect 8300 10310 8352 10362
rect 8364 10310 8416 10362
rect 8428 10310 8480 10362
rect 15946 10310 15998 10362
rect 16010 10310 16062 10362
rect 16074 10310 16126 10362
rect 16138 10310 16190 10362
rect 16202 10310 16254 10362
rect 23720 10310 23772 10362
rect 23784 10310 23836 10362
rect 23848 10310 23900 10362
rect 23912 10310 23964 10362
rect 23976 10310 24028 10362
rect 31494 10310 31546 10362
rect 31558 10310 31610 10362
rect 31622 10310 31674 10362
rect 31686 10310 31738 10362
rect 31750 10310 31802 10362
rect 4285 9766 4337 9818
rect 4349 9766 4401 9818
rect 4413 9766 4465 9818
rect 4477 9766 4529 9818
rect 4541 9766 4593 9818
rect 12059 9766 12111 9818
rect 12123 9766 12175 9818
rect 12187 9766 12239 9818
rect 12251 9766 12303 9818
rect 12315 9766 12367 9818
rect 19833 9766 19885 9818
rect 19897 9766 19949 9818
rect 19961 9766 20013 9818
rect 20025 9766 20077 9818
rect 20089 9766 20141 9818
rect 27607 9766 27659 9818
rect 27671 9766 27723 9818
rect 27735 9766 27787 9818
rect 27799 9766 27851 9818
rect 27863 9766 27915 9818
rect 8172 9222 8224 9274
rect 8236 9222 8288 9274
rect 8300 9222 8352 9274
rect 8364 9222 8416 9274
rect 8428 9222 8480 9274
rect 15946 9222 15998 9274
rect 16010 9222 16062 9274
rect 16074 9222 16126 9274
rect 16138 9222 16190 9274
rect 16202 9222 16254 9274
rect 23720 9222 23772 9274
rect 23784 9222 23836 9274
rect 23848 9222 23900 9274
rect 23912 9222 23964 9274
rect 23976 9222 24028 9274
rect 31494 9222 31546 9274
rect 31558 9222 31610 9274
rect 31622 9222 31674 9274
rect 31686 9222 31738 9274
rect 31750 9222 31802 9274
rect 4285 8678 4337 8730
rect 4349 8678 4401 8730
rect 4413 8678 4465 8730
rect 4477 8678 4529 8730
rect 4541 8678 4593 8730
rect 12059 8678 12111 8730
rect 12123 8678 12175 8730
rect 12187 8678 12239 8730
rect 12251 8678 12303 8730
rect 12315 8678 12367 8730
rect 19833 8678 19885 8730
rect 19897 8678 19949 8730
rect 19961 8678 20013 8730
rect 20025 8678 20077 8730
rect 20089 8678 20141 8730
rect 27607 8678 27659 8730
rect 27671 8678 27723 8730
rect 27735 8678 27787 8730
rect 27799 8678 27851 8730
rect 27863 8678 27915 8730
rect 8172 8134 8224 8186
rect 8236 8134 8288 8186
rect 8300 8134 8352 8186
rect 8364 8134 8416 8186
rect 8428 8134 8480 8186
rect 15946 8134 15998 8186
rect 16010 8134 16062 8186
rect 16074 8134 16126 8186
rect 16138 8134 16190 8186
rect 16202 8134 16254 8186
rect 23720 8134 23772 8186
rect 23784 8134 23836 8186
rect 23848 8134 23900 8186
rect 23912 8134 23964 8186
rect 23976 8134 24028 8186
rect 31494 8134 31546 8186
rect 31558 8134 31610 8186
rect 31622 8134 31674 8186
rect 31686 8134 31738 8186
rect 31750 8134 31802 8186
rect 4285 7590 4337 7642
rect 4349 7590 4401 7642
rect 4413 7590 4465 7642
rect 4477 7590 4529 7642
rect 4541 7590 4593 7642
rect 12059 7590 12111 7642
rect 12123 7590 12175 7642
rect 12187 7590 12239 7642
rect 12251 7590 12303 7642
rect 12315 7590 12367 7642
rect 19833 7590 19885 7642
rect 19897 7590 19949 7642
rect 19961 7590 20013 7642
rect 20025 7590 20077 7642
rect 20089 7590 20141 7642
rect 27607 7590 27659 7642
rect 27671 7590 27723 7642
rect 27735 7590 27787 7642
rect 27799 7590 27851 7642
rect 27863 7590 27915 7642
rect 8172 7046 8224 7098
rect 8236 7046 8288 7098
rect 8300 7046 8352 7098
rect 8364 7046 8416 7098
rect 8428 7046 8480 7098
rect 15946 7046 15998 7098
rect 16010 7046 16062 7098
rect 16074 7046 16126 7098
rect 16138 7046 16190 7098
rect 16202 7046 16254 7098
rect 23720 7046 23772 7098
rect 23784 7046 23836 7098
rect 23848 7046 23900 7098
rect 23912 7046 23964 7098
rect 23976 7046 24028 7098
rect 31494 7046 31546 7098
rect 31558 7046 31610 7098
rect 31622 7046 31674 7098
rect 31686 7046 31738 7098
rect 31750 7046 31802 7098
rect 4285 6502 4337 6554
rect 4349 6502 4401 6554
rect 4413 6502 4465 6554
rect 4477 6502 4529 6554
rect 4541 6502 4593 6554
rect 12059 6502 12111 6554
rect 12123 6502 12175 6554
rect 12187 6502 12239 6554
rect 12251 6502 12303 6554
rect 12315 6502 12367 6554
rect 19833 6502 19885 6554
rect 19897 6502 19949 6554
rect 19961 6502 20013 6554
rect 20025 6502 20077 6554
rect 20089 6502 20141 6554
rect 27607 6502 27659 6554
rect 27671 6502 27723 6554
rect 27735 6502 27787 6554
rect 27799 6502 27851 6554
rect 27863 6502 27915 6554
rect 8172 5958 8224 6010
rect 8236 5958 8288 6010
rect 8300 5958 8352 6010
rect 8364 5958 8416 6010
rect 8428 5958 8480 6010
rect 15946 5958 15998 6010
rect 16010 5958 16062 6010
rect 16074 5958 16126 6010
rect 16138 5958 16190 6010
rect 16202 5958 16254 6010
rect 23720 5958 23772 6010
rect 23784 5958 23836 6010
rect 23848 5958 23900 6010
rect 23912 5958 23964 6010
rect 23976 5958 24028 6010
rect 31494 5958 31546 6010
rect 31558 5958 31610 6010
rect 31622 5958 31674 6010
rect 31686 5958 31738 6010
rect 31750 5958 31802 6010
rect 4285 5414 4337 5466
rect 4349 5414 4401 5466
rect 4413 5414 4465 5466
rect 4477 5414 4529 5466
rect 4541 5414 4593 5466
rect 12059 5414 12111 5466
rect 12123 5414 12175 5466
rect 12187 5414 12239 5466
rect 12251 5414 12303 5466
rect 12315 5414 12367 5466
rect 19833 5414 19885 5466
rect 19897 5414 19949 5466
rect 19961 5414 20013 5466
rect 20025 5414 20077 5466
rect 20089 5414 20141 5466
rect 27607 5414 27659 5466
rect 27671 5414 27723 5466
rect 27735 5414 27787 5466
rect 27799 5414 27851 5466
rect 27863 5414 27915 5466
rect 8172 4870 8224 4922
rect 8236 4870 8288 4922
rect 8300 4870 8352 4922
rect 8364 4870 8416 4922
rect 8428 4870 8480 4922
rect 15946 4870 15998 4922
rect 16010 4870 16062 4922
rect 16074 4870 16126 4922
rect 16138 4870 16190 4922
rect 16202 4870 16254 4922
rect 23720 4870 23772 4922
rect 23784 4870 23836 4922
rect 23848 4870 23900 4922
rect 23912 4870 23964 4922
rect 23976 4870 24028 4922
rect 31494 4870 31546 4922
rect 31558 4870 31610 4922
rect 31622 4870 31674 4922
rect 31686 4870 31738 4922
rect 31750 4870 31802 4922
rect 4285 4326 4337 4378
rect 4349 4326 4401 4378
rect 4413 4326 4465 4378
rect 4477 4326 4529 4378
rect 4541 4326 4593 4378
rect 12059 4326 12111 4378
rect 12123 4326 12175 4378
rect 12187 4326 12239 4378
rect 12251 4326 12303 4378
rect 12315 4326 12367 4378
rect 19833 4326 19885 4378
rect 19897 4326 19949 4378
rect 19961 4326 20013 4378
rect 20025 4326 20077 4378
rect 20089 4326 20141 4378
rect 27607 4326 27659 4378
rect 27671 4326 27723 4378
rect 27735 4326 27787 4378
rect 27799 4326 27851 4378
rect 27863 4326 27915 4378
rect 8172 3782 8224 3834
rect 8236 3782 8288 3834
rect 8300 3782 8352 3834
rect 8364 3782 8416 3834
rect 8428 3782 8480 3834
rect 15946 3782 15998 3834
rect 16010 3782 16062 3834
rect 16074 3782 16126 3834
rect 16138 3782 16190 3834
rect 16202 3782 16254 3834
rect 23720 3782 23772 3834
rect 23784 3782 23836 3834
rect 23848 3782 23900 3834
rect 23912 3782 23964 3834
rect 23976 3782 24028 3834
rect 31494 3782 31546 3834
rect 31558 3782 31610 3834
rect 31622 3782 31674 3834
rect 31686 3782 31738 3834
rect 31750 3782 31802 3834
rect 4285 3238 4337 3290
rect 4349 3238 4401 3290
rect 4413 3238 4465 3290
rect 4477 3238 4529 3290
rect 4541 3238 4593 3290
rect 12059 3238 12111 3290
rect 12123 3238 12175 3290
rect 12187 3238 12239 3290
rect 12251 3238 12303 3290
rect 12315 3238 12367 3290
rect 19833 3238 19885 3290
rect 19897 3238 19949 3290
rect 19961 3238 20013 3290
rect 20025 3238 20077 3290
rect 20089 3238 20141 3290
rect 27607 3238 27659 3290
rect 27671 3238 27723 3290
rect 27735 3238 27787 3290
rect 27799 3238 27851 3290
rect 27863 3238 27915 3290
rect 8172 2694 8224 2746
rect 8236 2694 8288 2746
rect 8300 2694 8352 2746
rect 8364 2694 8416 2746
rect 8428 2694 8480 2746
rect 15946 2694 15998 2746
rect 16010 2694 16062 2746
rect 16074 2694 16126 2746
rect 16138 2694 16190 2746
rect 16202 2694 16254 2746
rect 23720 2694 23772 2746
rect 23784 2694 23836 2746
rect 23848 2694 23900 2746
rect 23912 2694 23964 2746
rect 23976 2694 24028 2746
rect 31494 2694 31546 2746
rect 31558 2694 31610 2746
rect 31622 2694 31674 2746
rect 31686 2694 31738 2746
rect 31750 2694 31802 2746
rect 4285 2150 4337 2202
rect 4349 2150 4401 2202
rect 4413 2150 4465 2202
rect 4477 2150 4529 2202
rect 4541 2150 4593 2202
rect 12059 2150 12111 2202
rect 12123 2150 12175 2202
rect 12187 2150 12239 2202
rect 12251 2150 12303 2202
rect 12315 2150 12367 2202
rect 19833 2150 19885 2202
rect 19897 2150 19949 2202
rect 19961 2150 20013 2202
rect 20025 2150 20077 2202
rect 20089 2150 20141 2202
rect 27607 2150 27659 2202
rect 27671 2150 27723 2202
rect 27735 2150 27787 2202
rect 27799 2150 27851 2202
rect 27863 2150 27915 2202
rect 8172 1606 8224 1658
rect 8236 1606 8288 1658
rect 8300 1606 8352 1658
rect 8364 1606 8416 1658
rect 8428 1606 8480 1658
rect 15946 1606 15998 1658
rect 16010 1606 16062 1658
rect 16074 1606 16126 1658
rect 16138 1606 16190 1658
rect 16202 1606 16254 1658
rect 23720 1606 23772 1658
rect 23784 1606 23836 1658
rect 23848 1606 23900 1658
rect 23912 1606 23964 1658
rect 23976 1606 24028 1658
rect 31494 1606 31546 1658
rect 31558 1606 31610 1658
rect 31622 1606 31674 1658
rect 31686 1606 31738 1658
rect 31750 1606 31802 1658
rect 4285 1062 4337 1114
rect 4349 1062 4401 1114
rect 4413 1062 4465 1114
rect 4477 1062 4529 1114
rect 4541 1062 4593 1114
rect 12059 1062 12111 1114
rect 12123 1062 12175 1114
rect 12187 1062 12239 1114
rect 12251 1062 12303 1114
rect 12315 1062 12367 1114
rect 19833 1062 19885 1114
rect 19897 1062 19949 1114
rect 19961 1062 20013 1114
rect 20025 1062 20077 1114
rect 20089 1062 20141 1114
rect 27607 1062 27659 1114
rect 27671 1062 27723 1114
rect 27735 1062 27787 1114
rect 27799 1062 27851 1114
rect 27863 1062 27915 1114
rect 8172 518 8224 570
rect 8236 518 8288 570
rect 8300 518 8352 570
rect 8364 518 8416 570
rect 8428 518 8480 570
rect 15946 518 15998 570
rect 16010 518 16062 570
rect 16074 518 16126 570
rect 16138 518 16190 570
rect 16202 518 16254 570
rect 23720 518 23772 570
rect 23784 518 23836 570
rect 23848 518 23900 570
rect 23912 518 23964 570
rect 23976 518 24028 570
rect 31494 518 31546 570
rect 31558 518 31610 570
rect 31622 518 31674 570
rect 31686 518 31738 570
rect 31750 518 31802 570
<< metal2 >>
rect 29182 22264 29238 22273
rect 29182 22199 29238 22208
rect 4526 21992 4582 22001
rect 8390 21992 8446 22001
rect 4582 21950 4660 21978
rect 4526 21927 4582 21936
rect 846 21856 902 21865
rect 846 21791 902 21800
rect 1582 21856 1638 21865
rect 1582 21791 1638 21800
rect 2318 21856 2374 21865
rect 2318 21791 2374 21800
rect 3238 21856 3294 21865
rect 3238 21791 3294 21800
rect 3790 21856 3846 21865
rect 3790 21791 3846 21800
rect 860 21690 888 21791
rect 1596 21690 1624 21791
rect 2332 21690 2360 21791
rect 3252 21690 3280 21791
rect 3804 21690 3832 21791
rect 4285 21788 4593 21797
rect 4285 21786 4291 21788
rect 4347 21786 4371 21788
rect 4427 21786 4451 21788
rect 4507 21786 4531 21788
rect 4587 21786 4593 21788
rect 4347 21734 4349 21786
rect 4529 21734 4531 21786
rect 4285 21732 4291 21734
rect 4347 21732 4371 21734
rect 4427 21732 4451 21734
rect 4507 21732 4531 21734
rect 4587 21732 4593 21734
rect 4285 21723 4593 21732
rect 4632 21690 4660 21950
rect 8390 21927 8446 21936
rect 16302 21992 16358 22001
rect 16302 21927 16358 21936
rect 27160 21956 27212 21962
rect 5262 21856 5318 21865
rect 5262 21791 5318 21800
rect 5998 21856 6054 21865
rect 5998 21791 6054 21800
rect 6734 21856 6790 21865
rect 6734 21791 6790 21800
rect 7470 21856 7526 21865
rect 7470 21791 7526 21800
rect 5276 21690 5304 21791
rect 6012 21690 6040 21791
rect 6748 21690 6776 21791
rect 7484 21690 7512 21791
rect 8404 21690 8432 21927
rect 8942 21856 8998 21865
rect 8942 21791 8998 21800
rect 9678 21856 9734 21865
rect 9678 21791 9734 21800
rect 10414 21856 10470 21865
rect 10414 21791 10470 21800
rect 11150 21856 11206 21865
rect 11150 21791 11206 21800
rect 11886 21856 11942 21865
rect 11886 21791 11942 21800
rect 12622 21856 12678 21865
rect 8956 21690 8984 21791
rect 9692 21690 9720 21791
rect 10428 21690 10456 21791
rect 11164 21690 11192 21791
rect 11900 21690 11928 21791
rect 12059 21788 12367 21797
rect 12622 21791 12678 21800
rect 13542 21856 13598 21865
rect 13542 21791 13598 21800
rect 14094 21856 14150 21865
rect 14094 21791 14150 21800
rect 14830 21856 14886 21865
rect 14830 21791 14886 21800
rect 15566 21856 15622 21865
rect 15566 21791 15622 21800
rect 12059 21786 12065 21788
rect 12121 21786 12145 21788
rect 12201 21786 12225 21788
rect 12281 21786 12305 21788
rect 12361 21786 12367 21788
rect 12121 21734 12123 21786
rect 12303 21734 12305 21786
rect 12059 21732 12065 21734
rect 12121 21732 12145 21734
rect 12201 21732 12225 21734
rect 12281 21732 12305 21734
rect 12361 21732 12367 21734
rect 12059 21723 12367 21732
rect 12636 21690 12664 21791
rect 13556 21690 13584 21791
rect 14108 21690 14136 21791
rect 14844 21690 14872 21791
rect 15580 21690 15608 21791
rect 16316 21690 16344 21927
rect 27160 21898 27212 21904
rect 29000 21956 29052 21962
rect 29000 21898 29052 21904
rect 26976 21888 27028 21894
rect 17038 21856 17094 21865
rect 26976 21830 27028 21836
rect 17038 21791 17094 21800
rect 17052 21690 17080 21791
rect 19833 21788 20141 21797
rect 19833 21786 19839 21788
rect 19895 21786 19919 21788
rect 19975 21786 19999 21788
rect 20055 21786 20079 21788
rect 20135 21786 20141 21788
rect 19895 21734 19897 21786
rect 20077 21734 20079 21786
rect 19833 21732 19839 21734
rect 19895 21732 19919 21734
rect 19975 21732 19999 21734
rect 20055 21732 20079 21734
rect 20135 21732 20141 21734
rect 19833 21723 20141 21732
rect 848 21684 900 21690
rect 848 21626 900 21632
rect 1584 21684 1636 21690
rect 1584 21626 1636 21632
rect 2320 21684 2372 21690
rect 2320 21626 2372 21632
rect 3240 21684 3292 21690
rect 3240 21626 3292 21632
rect 3792 21684 3844 21690
rect 3792 21626 3844 21632
rect 4620 21684 4672 21690
rect 4620 21626 4672 21632
rect 5264 21684 5316 21690
rect 5264 21626 5316 21632
rect 6000 21684 6052 21690
rect 6000 21626 6052 21632
rect 6736 21684 6788 21690
rect 6736 21626 6788 21632
rect 7472 21684 7524 21690
rect 7472 21626 7524 21632
rect 8392 21684 8444 21690
rect 8392 21626 8444 21632
rect 8944 21684 8996 21690
rect 8944 21626 8996 21632
rect 9680 21684 9732 21690
rect 9680 21626 9732 21632
rect 10416 21684 10468 21690
rect 10416 21626 10468 21632
rect 11152 21684 11204 21690
rect 11152 21626 11204 21632
rect 11888 21684 11940 21690
rect 11888 21626 11940 21632
rect 12624 21684 12676 21690
rect 12624 21626 12676 21632
rect 13544 21684 13596 21690
rect 13544 21626 13596 21632
rect 14096 21684 14148 21690
rect 14096 21626 14148 21632
rect 14832 21684 14884 21690
rect 14832 21626 14884 21632
rect 15568 21684 15620 21690
rect 15568 21626 15620 21632
rect 16304 21684 16356 21690
rect 16304 21626 16356 21632
rect 17040 21684 17092 21690
rect 17040 21626 17092 21632
rect 26988 21486 27016 21830
rect 27172 21554 27200 21898
rect 27607 21788 27915 21797
rect 27607 21786 27613 21788
rect 27669 21786 27693 21788
rect 27749 21786 27773 21788
rect 27829 21786 27853 21788
rect 27909 21786 27915 21788
rect 27669 21734 27671 21786
rect 27851 21734 27853 21786
rect 27607 21732 27613 21734
rect 27669 21732 27693 21734
rect 27749 21732 27773 21734
rect 27829 21732 27853 21734
rect 27909 21732 27915 21734
rect 27607 21723 27915 21732
rect 29012 21690 29040 21898
rect 29000 21684 29052 21690
rect 29000 21626 29052 21632
rect 27160 21548 27212 21554
rect 27160 21490 27212 21496
rect 29196 21486 29224 22199
rect 29552 21888 29604 21894
rect 29552 21830 29604 21836
rect 29734 21856 29790 21865
rect 29564 21690 29592 21830
rect 29734 21791 29790 21800
rect 29552 21684 29604 21690
rect 29552 21626 29604 21632
rect 29748 21486 29776 21791
rect 26976 21480 27028 21486
rect 26976 21422 27028 21428
rect 29184 21480 29236 21486
rect 29184 21422 29236 21428
rect 29736 21480 29788 21486
rect 29736 21422 29788 21428
rect 25688 21344 25740 21350
rect 25688 21286 25740 21292
rect 8172 21244 8480 21253
rect 8172 21242 8178 21244
rect 8234 21242 8258 21244
rect 8314 21242 8338 21244
rect 8394 21242 8418 21244
rect 8474 21242 8480 21244
rect 8234 21190 8236 21242
rect 8416 21190 8418 21242
rect 8172 21188 8178 21190
rect 8234 21188 8258 21190
rect 8314 21188 8338 21190
rect 8394 21188 8418 21190
rect 8474 21188 8480 21190
rect 8172 21179 8480 21188
rect 15946 21244 16254 21253
rect 15946 21242 15952 21244
rect 16008 21242 16032 21244
rect 16088 21242 16112 21244
rect 16168 21242 16192 21244
rect 16248 21242 16254 21244
rect 16008 21190 16010 21242
rect 16190 21190 16192 21242
rect 15946 21188 15952 21190
rect 16008 21188 16032 21190
rect 16088 21188 16112 21190
rect 16168 21188 16192 21190
rect 16248 21188 16254 21190
rect 15946 21179 16254 21188
rect 23720 21244 24028 21253
rect 23720 21242 23726 21244
rect 23782 21242 23806 21244
rect 23862 21242 23886 21244
rect 23942 21242 23966 21244
rect 24022 21242 24028 21244
rect 23782 21190 23784 21242
rect 23964 21190 23966 21242
rect 23720 21188 23726 21190
rect 23782 21188 23806 21190
rect 23862 21188 23886 21190
rect 23942 21188 23966 21190
rect 24022 21188 24028 21190
rect 23720 21179 24028 21188
rect 4285 20700 4593 20709
rect 4285 20698 4291 20700
rect 4347 20698 4371 20700
rect 4427 20698 4451 20700
rect 4507 20698 4531 20700
rect 4587 20698 4593 20700
rect 4347 20646 4349 20698
rect 4529 20646 4531 20698
rect 4285 20644 4291 20646
rect 4347 20644 4371 20646
rect 4427 20644 4451 20646
rect 4507 20644 4531 20646
rect 4587 20644 4593 20646
rect 4285 20635 4593 20644
rect 12059 20700 12367 20709
rect 12059 20698 12065 20700
rect 12121 20698 12145 20700
rect 12201 20698 12225 20700
rect 12281 20698 12305 20700
rect 12361 20698 12367 20700
rect 12121 20646 12123 20698
rect 12303 20646 12305 20698
rect 12059 20644 12065 20646
rect 12121 20644 12145 20646
rect 12201 20644 12225 20646
rect 12281 20644 12305 20646
rect 12361 20644 12367 20646
rect 12059 20635 12367 20644
rect 19833 20700 20141 20709
rect 19833 20698 19839 20700
rect 19895 20698 19919 20700
rect 19975 20698 19999 20700
rect 20055 20698 20079 20700
rect 20135 20698 20141 20700
rect 19895 20646 19897 20698
rect 20077 20646 20079 20698
rect 19833 20644 19839 20646
rect 19895 20644 19919 20646
rect 19975 20644 19999 20646
rect 20055 20644 20079 20646
rect 20135 20644 20141 20646
rect 19833 20635 20141 20644
rect 8172 20156 8480 20165
rect 8172 20154 8178 20156
rect 8234 20154 8258 20156
rect 8314 20154 8338 20156
rect 8394 20154 8418 20156
rect 8474 20154 8480 20156
rect 8234 20102 8236 20154
rect 8416 20102 8418 20154
rect 8172 20100 8178 20102
rect 8234 20100 8258 20102
rect 8314 20100 8338 20102
rect 8394 20100 8418 20102
rect 8474 20100 8480 20102
rect 8172 20091 8480 20100
rect 15946 20156 16254 20165
rect 15946 20154 15952 20156
rect 16008 20154 16032 20156
rect 16088 20154 16112 20156
rect 16168 20154 16192 20156
rect 16248 20154 16254 20156
rect 16008 20102 16010 20154
rect 16190 20102 16192 20154
rect 15946 20100 15952 20102
rect 16008 20100 16032 20102
rect 16088 20100 16112 20102
rect 16168 20100 16192 20102
rect 16248 20100 16254 20102
rect 15946 20091 16254 20100
rect 23720 20156 24028 20165
rect 23720 20154 23726 20156
rect 23782 20154 23806 20156
rect 23862 20154 23886 20156
rect 23942 20154 23966 20156
rect 24022 20154 24028 20156
rect 23782 20102 23784 20154
rect 23964 20102 23966 20154
rect 23720 20100 23726 20102
rect 23782 20100 23806 20102
rect 23862 20100 23886 20102
rect 23942 20100 23966 20102
rect 24022 20100 24028 20102
rect 23720 20091 24028 20100
rect 4285 19612 4593 19621
rect 4285 19610 4291 19612
rect 4347 19610 4371 19612
rect 4427 19610 4451 19612
rect 4507 19610 4531 19612
rect 4587 19610 4593 19612
rect 4347 19558 4349 19610
rect 4529 19558 4531 19610
rect 4285 19556 4291 19558
rect 4347 19556 4371 19558
rect 4427 19556 4451 19558
rect 4507 19556 4531 19558
rect 4587 19556 4593 19558
rect 4285 19547 4593 19556
rect 12059 19612 12367 19621
rect 12059 19610 12065 19612
rect 12121 19610 12145 19612
rect 12201 19610 12225 19612
rect 12281 19610 12305 19612
rect 12361 19610 12367 19612
rect 12121 19558 12123 19610
rect 12303 19558 12305 19610
rect 12059 19556 12065 19558
rect 12121 19556 12145 19558
rect 12201 19556 12225 19558
rect 12281 19556 12305 19558
rect 12361 19556 12367 19558
rect 12059 19547 12367 19556
rect 19833 19612 20141 19621
rect 19833 19610 19839 19612
rect 19895 19610 19919 19612
rect 19975 19610 19999 19612
rect 20055 19610 20079 19612
rect 20135 19610 20141 19612
rect 19895 19558 19897 19610
rect 20077 19558 20079 19610
rect 19833 19556 19839 19558
rect 19895 19556 19919 19558
rect 19975 19556 19999 19558
rect 20055 19556 20079 19558
rect 20135 19556 20141 19558
rect 19833 19547 20141 19556
rect 25700 19281 25728 21286
rect 31494 21244 31802 21253
rect 31494 21242 31500 21244
rect 31556 21242 31580 21244
rect 31636 21242 31660 21244
rect 31716 21242 31740 21244
rect 31796 21242 31802 21244
rect 31556 21190 31558 21242
rect 31738 21190 31740 21242
rect 31494 21188 31500 21190
rect 31556 21188 31580 21190
rect 31636 21188 31660 21190
rect 31716 21188 31740 21190
rect 31796 21188 31802 21190
rect 31494 21179 31802 21188
rect 27607 20700 27915 20709
rect 27607 20698 27613 20700
rect 27669 20698 27693 20700
rect 27749 20698 27773 20700
rect 27829 20698 27853 20700
rect 27909 20698 27915 20700
rect 27669 20646 27671 20698
rect 27851 20646 27853 20698
rect 27607 20644 27613 20646
rect 27669 20644 27693 20646
rect 27749 20644 27773 20646
rect 27829 20644 27853 20646
rect 27909 20644 27915 20646
rect 27607 20635 27915 20644
rect 31494 20156 31802 20165
rect 31494 20154 31500 20156
rect 31556 20154 31580 20156
rect 31636 20154 31660 20156
rect 31716 20154 31740 20156
rect 31796 20154 31802 20156
rect 31556 20102 31558 20154
rect 31738 20102 31740 20154
rect 31494 20100 31500 20102
rect 31556 20100 31580 20102
rect 31636 20100 31660 20102
rect 31716 20100 31740 20102
rect 31796 20100 31802 20102
rect 31494 20091 31802 20100
rect 27607 19612 27915 19621
rect 27607 19610 27613 19612
rect 27669 19610 27693 19612
rect 27749 19610 27773 19612
rect 27829 19610 27853 19612
rect 27909 19610 27915 19612
rect 27669 19558 27671 19610
rect 27851 19558 27853 19610
rect 27607 19556 27613 19558
rect 27669 19556 27693 19558
rect 27749 19556 27773 19558
rect 27829 19556 27853 19558
rect 27909 19556 27915 19558
rect 27607 19547 27915 19556
rect 25686 19272 25742 19281
rect 25686 19207 25742 19216
rect 8172 19068 8480 19077
rect 8172 19066 8178 19068
rect 8234 19066 8258 19068
rect 8314 19066 8338 19068
rect 8394 19066 8418 19068
rect 8474 19066 8480 19068
rect 8234 19014 8236 19066
rect 8416 19014 8418 19066
rect 8172 19012 8178 19014
rect 8234 19012 8258 19014
rect 8314 19012 8338 19014
rect 8394 19012 8418 19014
rect 8474 19012 8480 19014
rect 8172 19003 8480 19012
rect 15946 19068 16254 19077
rect 15946 19066 15952 19068
rect 16008 19066 16032 19068
rect 16088 19066 16112 19068
rect 16168 19066 16192 19068
rect 16248 19066 16254 19068
rect 16008 19014 16010 19066
rect 16190 19014 16192 19066
rect 15946 19012 15952 19014
rect 16008 19012 16032 19014
rect 16088 19012 16112 19014
rect 16168 19012 16192 19014
rect 16248 19012 16254 19014
rect 15946 19003 16254 19012
rect 23720 19068 24028 19077
rect 23720 19066 23726 19068
rect 23782 19066 23806 19068
rect 23862 19066 23886 19068
rect 23942 19066 23966 19068
rect 24022 19066 24028 19068
rect 23782 19014 23784 19066
rect 23964 19014 23966 19066
rect 23720 19012 23726 19014
rect 23782 19012 23806 19014
rect 23862 19012 23886 19014
rect 23942 19012 23966 19014
rect 24022 19012 24028 19014
rect 23720 19003 24028 19012
rect 31494 19068 31802 19077
rect 31494 19066 31500 19068
rect 31556 19066 31580 19068
rect 31636 19066 31660 19068
rect 31716 19066 31740 19068
rect 31796 19066 31802 19068
rect 31556 19014 31558 19066
rect 31738 19014 31740 19066
rect 31494 19012 31500 19014
rect 31556 19012 31580 19014
rect 31636 19012 31660 19014
rect 31716 19012 31740 19014
rect 31796 19012 31802 19014
rect 31494 19003 31802 19012
rect 4285 18524 4593 18533
rect 4285 18522 4291 18524
rect 4347 18522 4371 18524
rect 4427 18522 4451 18524
rect 4507 18522 4531 18524
rect 4587 18522 4593 18524
rect 4347 18470 4349 18522
rect 4529 18470 4531 18522
rect 4285 18468 4291 18470
rect 4347 18468 4371 18470
rect 4427 18468 4451 18470
rect 4507 18468 4531 18470
rect 4587 18468 4593 18470
rect 4285 18459 4593 18468
rect 12059 18524 12367 18533
rect 12059 18522 12065 18524
rect 12121 18522 12145 18524
rect 12201 18522 12225 18524
rect 12281 18522 12305 18524
rect 12361 18522 12367 18524
rect 12121 18470 12123 18522
rect 12303 18470 12305 18522
rect 12059 18468 12065 18470
rect 12121 18468 12145 18470
rect 12201 18468 12225 18470
rect 12281 18468 12305 18470
rect 12361 18468 12367 18470
rect 12059 18459 12367 18468
rect 19833 18524 20141 18533
rect 19833 18522 19839 18524
rect 19895 18522 19919 18524
rect 19975 18522 19999 18524
rect 20055 18522 20079 18524
rect 20135 18522 20141 18524
rect 19895 18470 19897 18522
rect 20077 18470 20079 18522
rect 19833 18468 19839 18470
rect 19895 18468 19919 18470
rect 19975 18468 19999 18470
rect 20055 18468 20079 18470
rect 20135 18468 20141 18470
rect 19833 18459 20141 18468
rect 27607 18524 27915 18533
rect 27607 18522 27613 18524
rect 27669 18522 27693 18524
rect 27749 18522 27773 18524
rect 27829 18522 27853 18524
rect 27909 18522 27915 18524
rect 27669 18470 27671 18522
rect 27851 18470 27853 18522
rect 27607 18468 27613 18470
rect 27669 18468 27693 18470
rect 27749 18468 27773 18470
rect 27829 18468 27853 18470
rect 27909 18468 27915 18470
rect 27607 18459 27915 18468
rect 8172 17980 8480 17989
rect 8172 17978 8178 17980
rect 8234 17978 8258 17980
rect 8314 17978 8338 17980
rect 8394 17978 8418 17980
rect 8474 17978 8480 17980
rect 8234 17926 8236 17978
rect 8416 17926 8418 17978
rect 8172 17924 8178 17926
rect 8234 17924 8258 17926
rect 8314 17924 8338 17926
rect 8394 17924 8418 17926
rect 8474 17924 8480 17926
rect 8172 17915 8480 17924
rect 15946 17980 16254 17989
rect 15946 17978 15952 17980
rect 16008 17978 16032 17980
rect 16088 17978 16112 17980
rect 16168 17978 16192 17980
rect 16248 17978 16254 17980
rect 16008 17926 16010 17978
rect 16190 17926 16192 17978
rect 15946 17924 15952 17926
rect 16008 17924 16032 17926
rect 16088 17924 16112 17926
rect 16168 17924 16192 17926
rect 16248 17924 16254 17926
rect 15946 17915 16254 17924
rect 23720 17980 24028 17989
rect 23720 17978 23726 17980
rect 23782 17978 23806 17980
rect 23862 17978 23886 17980
rect 23942 17978 23966 17980
rect 24022 17978 24028 17980
rect 23782 17926 23784 17978
rect 23964 17926 23966 17978
rect 23720 17924 23726 17926
rect 23782 17924 23806 17926
rect 23862 17924 23886 17926
rect 23942 17924 23966 17926
rect 24022 17924 24028 17926
rect 23720 17915 24028 17924
rect 31494 17980 31802 17989
rect 31494 17978 31500 17980
rect 31556 17978 31580 17980
rect 31636 17978 31660 17980
rect 31716 17978 31740 17980
rect 31796 17978 31802 17980
rect 31556 17926 31558 17978
rect 31738 17926 31740 17978
rect 31494 17924 31500 17926
rect 31556 17924 31580 17926
rect 31636 17924 31660 17926
rect 31716 17924 31740 17926
rect 31796 17924 31802 17926
rect 31494 17915 31802 17924
rect 4285 17436 4593 17445
rect 4285 17434 4291 17436
rect 4347 17434 4371 17436
rect 4427 17434 4451 17436
rect 4507 17434 4531 17436
rect 4587 17434 4593 17436
rect 4347 17382 4349 17434
rect 4529 17382 4531 17434
rect 4285 17380 4291 17382
rect 4347 17380 4371 17382
rect 4427 17380 4451 17382
rect 4507 17380 4531 17382
rect 4587 17380 4593 17382
rect 4285 17371 4593 17380
rect 12059 17436 12367 17445
rect 12059 17434 12065 17436
rect 12121 17434 12145 17436
rect 12201 17434 12225 17436
rect 12281 17434 12305 17436
rect 12361 17434 12367 17436
rect 12121 17382 12123 17434
rect 12303 17382 12305 17434
rect 12059 17380 12065 17382
rect 12121 17380 12145 17382
rect 12201 17380 12225 17382
rect 12281 17380 12305 17382
rect 12361 17380 12367 17382
rect 12059 17371 12367 17380
rect 19833 17436 20141 17445
rect 19833 17434 19839 17436
rect 19895 17434 19919 17436
rect 19975 17434 19999 17436
rect 20055 17434 20079 17436
rect 20135 17434 20141 17436
rect 19895 17382 19897 17434
rect 20077 17382 20079 17434
rect 19833 17380 19839 17382
rect 19895 17380 19919 17382
rect 19975 17380 19999 17382
rect 20055 17380 20079 17382
rect 20135 17380 20141 17382
rect 19833 17371 20141 17380
rect 27607 17436 27915 17445
rect 27607 17434 27613 17436
rect 27669 17434 27693 17436
rect 27749 17434 27773 17436
rect 27829 17434 27853 17436
rect 27909 17434 27915 17436
rect 27669 17382 27671 17434
rect 27851 17382 27853 17434
rect 27607 17380 27613 17382
rect 27669 17380 27693 17382
rect 27749 17380 27773 17382
rect 27829 17380 27853 17382
rect 27909 17380 27915 17382
rect 27607 17371 27915 17380
rect 8172 16892 8480 16901
rect 8172 16890 8178 16892
rect 8234 16890 8258 16892
rect 8314 16890 8338 16892
rect 8394 16890 8418 16892
rect 8474 16890 8480 16892
rect 8234 16838 8236 16890
rect 8416 16838 8418 16890
rect 8172 16836 8178 16838
rect 8234 16836 8258 16838
rect 8314 16836 8338 16838
rect 8394 16836 8418 16838
rect 8474 16836 8480 16838
rect 8172 16827 8480 16836
rect 15946 16892 16254 16901
rect 15946 16890 15952 16892
rect 16008 16890 16032 16892
rect 16088 16890 16112 16892
rect 16168 16890 16192 16892
rect 16248 16890 16254 16892
rect 16008 16838 16010 16890
rect 16190 16838 16192 16890
rect 15946 16836 15952 16838
rect 16008 16836 16032 16838
rect 16088 16836 16112 16838
rect 16168 16836 16192 16838
rect 16248 16836 16254 16838
rect 15946 16827 16254 16836
rect 23720 16892 24028 16901
rect 23720 16890 23726 16892
rect 23782 16890 23806 16892
rect 23862 16890 23886 16892
rect 23942 16890 23966 16892
rect 24022 16890 24028 16892
rect 23782 16838 23784 16890
rect 23964 16838 23966 16890
rect 23720 16836 23726 16838
rect 23782 16836 23806 16838
rect 23862 16836 23886 16838
rect 23942 16836 23966 16838
rect 24022 16836 24028 16838
rect 23720 16827 24028 16836
rect 31494 16892 31802 16901
rect 31494 16890 31500 16892
rect 31556 16890 31580 16892
rect 31636 16890 31660 16892
rect 31716 16890 31740 16892
rect 31796 16890 31802 16892
rect 31556 16838 31558 16890
rect 31738 16838 31740 16890
rect 31494 16836 31500 16838
rect 31556 16836 31580 16838
rect 31636 16836 31660 16838
rect 31716 16836 31740 16838
rect 31796 16836 31802 16838
rect 31494 16827 31802 16836
rect 4285 16348 4593 16357
rect 4285 16346 4291 16348
rect 4347 16346 4371 16348
rect 4427 16346 4451 16348
rect 4507 16346 4531 16348
rect 4587 16346 4593 16348
rect 4347 16294 4349 16346
rect 4529 16294 4531 16346
rect 4285 16292 4291 16294
rect 4347 16292 4371 16294
rect 4427 16292 4451 16294
rect 4507 16292 4531 16294
rect 4587 16292 4593 16294
rect 4285 16283 4593 16292
rect 12059 16348 12367 16357
rect 12059 16346 12065 16348
rect 12121 16346 12145 16348
rect 12201 16346 12225 16348
rect 12281 16346 12305 16348
rect 12361 16346 12367 16348
rect 12121 16294 12123 16346
rect 12303 16294 12305 16346
rect 12059 16292 12065 16294
rect 12121 16292 12145 16294
rect 12201 16292 12225 16294
rect 12281 16292 12305 16294
rect 12361 16292 12367 16294
rect 12059 16283 12367 16292
rect 19833 16348 20141 16357
rect 19833 16346 19839 16348
rect 19895 16346 19919 16348
rect 19975 16346 19999 16348
rect 20055 16346 20079 16348
rect 20135 16346 20141 16348
rect 19895 16294 19897 16346
rect 20077 16294 20079 16346
rect 19833 16292 19839 16294
rect 19895 16292 19919 16294
rect 19975 16292 19999 16294
rect 20055 16292 20079 16294
rect 20135 16292 20141 16294
rect 19833 16283 20141 16292
rect 27607 16348 27915 16357
rect 27607 16346 27613 16348
rect 27669 16346 27693 16348
rect 27749 16346 27773 16348
rect 27829 16346 27853 16348
rect 27909 16346 27915 16348
rect 27669 16294 27671 16346
rect 27851 16294 27853 16346
rect 27607 16292 27613 16294
rect 27669 16292 27693 16294
rect 27749 16292 27773 16294
rect 27829 16292 27853 16294
rect 27909 16292 27915 16294
rect 27607 16283 27915 16292
rect 8172 15804 8480 15813
rect 8172 15802 8178 15804
rect 8234 15802 8258 15804
rect 8314 15802 8338 15804
rect 8394 15802 8418 15804
rect 8474 15802 8480 15804
rect 8234 15750 8236 15802
rect 8416 15750 8418 15802
rect 8172 15748 8178 15750
rect 8234 15748 8258 15750
rect 8314 15748 8338 15750
rect 8394 15748 8418 15750
rect 8474 15748 8480 15750
rect 8172 15739 8480 15748
rect 15946 15804 16254 15813
rect 15946 15802 15952 15804
rect 16008 15802 16032 15804
rect 16088 15802 16112 15804
rect 16168 15802 16192 15804
rect 16248 15802 16254 15804
rect 16008 15750 16010 15802
rect 16190 15750 16192 15802
rect 15946 15748 15952 15750
rect 16008 15748 16032 15750
rect 16088 15748 16112 15750
rect 16168 15748 16192 15750
rect 16248 15748 16254 15750
rect 15946 15739 16254 15748
rect 23720 15804 24028 15813
rect 23720 15802 23726 15804
rect 23782 15802 23806 15804
rect 23862 15802 23886 15804
rect 23942 15802 23966 15804
rect 24022 15802 24028 15804
rect 23782 15750 23784 15802
rect 23964 15750 23966 15802
rect 23720 15748 23726 15750
rect 23782 15748 23806 15750
rect 23862 15748 23886 15750
rect 23942 15748 23966 15750
rect 24022 15748 24028 15750
rect 23720 15739 24028 15748
rect 31494 15804 31802 15813
rect 31494 15802 31500 15804
rect 31556 15802 31580 15804
rect 31636 15802 31660 15804
rect 31716 15802 31740 15804
rect 31796 15802 31802 15804
rect 31556 15750 31558 15802
rect 31738 15750 31740 15802
rect 31494 15748 31500 15750
rect 31556 15748 31580 15750
rect 31636 15748 31660 15750
rect 31716 15748 31740 15750
rect 31796 15748 31802 15750
rect 31494 15739 31802 15748
rect 4285 15260 4593 15269
rect 4285 15258 4291 15260
rect 4347 15258 4371 15260
rect 4427 15258 4451 15260
rect 4507 15258 4531 15260
rect 4587 15258 4593 15260
rect 4347 15206 4349 15258
rect 4529 15206 4531 15258
rect 4285 15204 4291 15206
rect 4347 15204 4371 15206
rect 4427 15204 4451 15206
rect 4507 15204 4531 15206
rect 4587 15204 4593 15206
rect 4285 15195 4593 15204
rect 12059 15260 12367 15269
rect 12059 15258 12065 15260
rect 12121 15258 12145 15260
rect 12201 15258 12225 15260
rect 12281 15258 12305 15260
rect 12361 15258 12367 15260
rect 12121 15206 12123 15258
rect 12303 15206 12305 15258
rect 12059 15204 12065 15206
rect 12121 15204 12145 15206
rect 12201 15204 12225 15206
rect 12281 15204 12305 15206
rect 12361 15204 12367 15206
rect 12059 15195 12367 15204
rect 19833 15260 20141 15269
rect 19833 15258 19839 15260
rect 19895 15258 19919 15260
rect 19975 15258 19999 15260
rect 20055 15258 20079 15260
rect 20135 15258 20141 15260
rect 19895 15206 19897 15258
rect 20077 15206 20079 15258
rect 19833 15204 19839 15206
rect 19895 15204 19919 15206
rect 19975 15204 19999 15206
rect 20055 15204 20079 15206
rect 20135 15204 20141 15206
rect 19833 15195 20141 15204
rect 27607 15260 27915 15269
rect 27607 15258 27613 15260
rect 27669 15258 27693 15260
rect 27749 15258 27773 15260
rect 27829 15258 27853 15260
rect 27909 15258 27915 15260
rect 27669 15206 27671 15258
rect 27851 15206 27853 15258
rect 27607 15204 27613 15206
rect 27669 15204 27693 15206
rect 27749 15204 27773 15206
rect 27829 15204 27853 15206
rect 27909 15204 27915 15206
rect 27607 15195 27915 15204
rect 8172 14716 8480 14725
rect 8172 14714 8178 14716
rect 8234 14714 8258 14716
rect 8314 14714 8338 14716
rect 8394 14714 8418 14716
rect 8474 14714 8480 14716
rect 8234 14662 8236 14714
rect 8416 14662 8418 14714
rect 8172 14660 8178 14662
rect 8234 14660 8258 14662
rect 8314 14660 8338 14662
rect 8394 14660 8418 14662
rect 8474 14660 8480 14662
rect 8172 14651 8480 14660
rect 15946 14716 16254 14725
rect 15946 14714 15952 14716
rect 16008 14714 16032 14716
rect 16088 14714 16112 14716
rect 16168 14714 16192 14716
rect 16248 14714 16254 14716
rect 16008 14662 16010 14714
rect 16190 14662 16192 14714
rect 15946 14660 15952 14662
rect 16008 14660 16032 14662
rect 16088 14660 16112 14662
rect 16168 14660 16192 14662
rect 16248 14660 16254 14662
rect 15946 14651 16254 14660
rect 23720 14716 24028 14725
rect 23720 14714 23726 14716
rect 23782 14714 23806 14716
rect 23862 14714 23886 14716
rect 23942 14714 23966 14716
rect 24022 14714 24028 14716
rect 23782 14662 23784 14714
rect 23964 14662 23966 14714
rect 23720 14660 23726 14662
rect 23782 14660 23806 14662
rect 23862 14660 23886 14662
rect 23942 14660 23966 14662
rect 24022 14660 24028 14662
rect 23720 14651 24028 14660
rect 31494 14716 31802 14725
rect 31494 14714 31500 14716
rect 31556 14714 31580 14716
rect 31636 14714 31660 14716
rect 31716 14714 31740 14716
rect 31796 14714 31802 14716
rect 31556 14662 31558 14714
rect 31738 14662 31740 14714
rect 31494 14660 31500 14662
rect 31556 14660 31580 14662
rect 31636 14660 31660 14662
rect 31716 14660 31740 14662
rect 31796 14660 31802 14662
rect 31494 14651 31802 14660
rect 4285 14172 4593 14181
rect 4285 14170 4291 14172
rect 4347 14170 4371 14172
rect 4427 14170 4451 14172
rect 4507 14170 4531 14172
rect 4587 14170 4593 14172
rect 4347 14118 4349 14170
rect 4529 14118 4531 14170
rect 4285 14116 4291 14118
rect 4347 14116 4371 14118
rect 4427 14116 4451 14118
rect 4507 14116 4531 14118
rect 4587 14116 4593 14118
rect 4285 14107 4593 14116
rect 12059 14172 12367 14181
rect 12059 14170 12065 14172
rect 12121 14170 12145 14172
rect 12201 14170 12225 14172
rect 12281 14170 12305 14172
rect 12361 14170 12367 14172
rect 12121 14118 12123 14170
rect 12303 14118 12305 14170
rect 12059 14116 12065 14118
rect 12121 14116 12145 14118
rect 12201 14116 12225 14118
rect 12281 14116 12305 14118
rect 12361 14116 12367 14118
rect 12059 14107 12367 14116
rect 19833 14172 20141 14181
rect 19833 14170 19839 14172
rect 19895 14170 19919 14172
rect 19975 14170 19999 14172
rect 20055 14170 20079 14172
rect 20135 14170 20141 14172
rect 19895 14118 19897 14170
rect 20077 14118 20079 14170
rect 19833 14116 19839 14118
rect 19895 14116 19919 14118
rect 19975 14116 19999 14118
rect 20055 14116 20079 14118
rect 20135 14116 20141 14118
rect 19833 14107 20141 14116
rect 27607 14172 27915 14181
rect 27607 14170 27613 14172
rect 27669 14170 27693 14172
rect 27749 14170 27773 14172
rect 27829 14170 27853 14172
rect 27909 14170 27915 14172
rect 27669 14118 27671 14170
rect 27851 14118 27853 14170
rect 27607 14116 27613 14118
rect 27669 14116 27693 14118
rect 27749 14116 27773 14118
rect 27829 14116 27853 14118
rect 27909 14116 27915 14118
rect 27607 14107 27915 14116
rect 8172 13628 8480 13637
rect 8172 13626 8178 13628
rect 8234 13626 8258 13628
rect 8314 13626 8338 13628
rect 8394 13626 8418 13628
rect 8474 13626 8480 13628
rect 8234 13574 8236 13626
rect 8416 13574 8418 13626
rect 8172 13572 8178 13574
rect 8234 13572 8258 13574
rect 8314 13572 8338 13574
rect 8394 13572 8418 13574
rect 8474 13572 8480 13574
rect 8172 13563 8480 13572
rect 15946 13628 16254 13637
rect 15946 13626 15952 13628
rect 16008 13626 16032 13628
rect 16088 13626 16112 13628
rect 16168 13626 16192 13628
rect 16248 13626 16254 13628
rect 16008 13574 16010 13626
rect 16190 13574 16192 13626
rect 15946 13572 15952 13574
rect 16008 13572 16032 13574
rect 16088 13572 16112 13574
rect 16168 13572 16192 13574
rect 16248 13572 16254 13574
rect 15946 13563 16254 13572
rect 23720 13628 24028 13637
rect 23720 13626 23726 13628
rect 23782 13626 23806 13628
rect 23862 13626 23886 13628
rect 23942 13626 23966 13628
rect 24022 13626 24028 13628
rect 23782 13574 23784 13626
rect 23964 13574 23966 13626
rect 23720 13572 23726 13574
rect 23782 13572 23806 13574
rect 23862 13572 23886 13574
rect 23942 13572 23966 13574
rect 24022 13572 24028 13574
rect 23720 13563 24028 13572
rect 31494 13628 31802 13637
rect 31494 13626 31500 13628
rect 31556 13626 31580 13628
rect 31636 13626 31660 13628
rect 31716 13626 31740 13628
rect 31796 13626 31802 13628
rect 31556 13574 31558 13626
rect 31738 13574 31740 13626
rect 31494 13572 31500 13574
rect 31556 13572 31580 13574
rect 31636 13572 31660 13574
rect 31716 13572 31740 13574
rect 31796 13572 31802 13574
rect 31494 13563 31802 13572
rect 4285 13084 4593 13093
rect 4285 13082 4291 13084
rect 4347 13082 4371 13084
rect 4427 13082 4451 13084
rect 4507 13082 4531 13084
rect 4587 13082 4593 13084
rect 4347 13030 4349 13082
rect 4529 13030 4531 13082
rect 4285 13028 4291 13030
rect 4347 13028 4371 13030
rect 4427 13028 4451 13030
rect 4507 13028 4531 13030
rect 4587 13028 4593 13030
rect 4285 13019 4593 13028
rect 12059 13084 12367 13093
rect 12059 13082 12065 13084
rect 12121 13082 12145 13084
rect 12201 13082 12225 13084
rect 12281 13082 12305 13084
rect 12361 13082 12367 13084
rect 12121 13030 12123 13082
rect 12303 13030 12305 13082
rect 12059 13028 12065 13030
rect 12121 13028 12145 13030
rect 12201 13028 12225 13030
rect 12281 13028 12305 13030
rect 12361 13028 12367 13030
rect 12059 13019 12367 13028
rect 19833 13084 20141 13093
rect 19833 13082 19839 13084
rect 19895 13082 19919 13084
rect 19975 13082 19999 13084
rect 20055 13082 20079 13084
rect 20135 13082 20141 13084
rect 19895 13030 19897 13082
rect 20077 13030 20079 13082
rect 19833 13028 19839 13030
rect 19895 13028 19919 13030
rect 19975 13028 19999 13030
rect 20055 13028 20079 13030
rect 20135 13028 20141 13030
rect 19833 13019 20141 13028
rect 27607 13084 27915 13093
rect 27607 13082 27613 13084
rect 27669 13082 27693 13084
rect 27749 13082 27773 13084
rect 27829 13082 27853 13084
rect 27909 13082 27915 13084
rect 27669 13030 27671 13082
rect 27851 13030 27853 13082
rect 27607 13028 27613 13030
rect 27669 13028 27693 13030
rect 27749 13028 27773 13030
rect 27829 13028 27853 13030
rect 27909 13028 27915 13030
rect 27607 13019 27915 13028
rect 8172 12540 8480 12549
rect 8172 12538 8178 12540
rect 8234 12538 8258 12540
rect 8314 12538 8338 12540
rect 8394 12538 8418 12540
rect 8474 12538 8480 12540
rect 8234 12486 8236 12538
rect 8416 12486 8418 12538
rect 8172 12484 8178 12486
rect 8234 12484 8258 12486
rect 8314 12484 8338 12486
rect 8394 12484 8418 12486
rect 8474 12484 8480 12486
rect 8172 12475 8480 12484
rect 15946 12540 16254 12549
rect 15946 12538 15952 12540
rect 16008 12538 16032 12540
rect 16088 12538 16112 12540
rect 16168 12538 16192 12540
rect 16248 12538 16254 12540
rect 16008 12486 16010 12538
rect 16190 12486 16192 12538
rect 15946 12484 15952 12486
rect 16008 12484 16032 12486
rect 16088 12484 16112 12486
rect 16168 12484 16192 12486
rect 16248 12484 16254 12486
rect 15946 12475 16254 12484
rect 23720 12540 24028 12549
rect 23720 12538 23726 12540
rect 23782 12538 23806 12540
rect 23862 12538 23886 12540
rect 23942 12538 23966 12540
rect 24022 12538 24028 12540
rect 23782 12486 23784 12538
rect 23964 12486 23966 12538
rect 23720 12484 23726 12486
rect 23782 12484 23806 12486
rect 23862 12484 23886 12486
rect 23942 12484 23966 12486
rect 24022 12484 24028 12486
rect 23720 12475 24028 12484
rect 31494 12540 31802 12549
rect 31494 12538 31500 12540
rect 31556 12538 31580 12540
rect 31636 12538 31660 12540
rect 31716 12538 31740 12540
rect 31796 12538 31802 12540
rect 31556 12486 31558 12538
rect 31738 12486 31740 12538
rect 31494 12484 31500 12486
rect 31556 12484 31580 12486
rect 31636 12484 31660 12486
rect 31716 12484 31740 12486
rect 31796 12484 31802 12486
rect 31494 12475 31802 12484
rect 4285 11996 4593 12005
rect 4285 11994 4291 11996
rect 4347 11994 4371 11996
rect 4427 11994 4451 11996
rect 4507 11994 4531 11996
rect 4587 11994 4593 11996
rect 4347 11942 4349 11994
rect 4529 11942 4531 11994
rect 4285 11940 4291 11942
rect 4347 11940 4371 11942
rect 4427 11940 4451 11942
rect 4507 11940 4531 11942
rect 4587 11940 4593 11942
rect 4285 11931 4593 11940
rect 12059 11996 12367 12005
rect 12059 11994 12065 11996
rect 12121 11994 12145 11996
rect 12201 11994 12225 11996
rect 12281 11994 12305 11996
rect 12361 11994 12367 11996
rect 12121 11942 12123 11994
rect 12303 11942 12305 11994
rect 12059 11940 12065 11942
rect 12121 11940 12145 11942
rect 12201 11940 12225 11942
rect 12281 11940 12305 11942
rect 12361 11940 12367 11942
rect 12059 11931 12367 11940
rect 19833 11996 20141 12005
rect 19833 11994 19839 11996
rect 19895 11994 19919 11996
rect 19975 11994 19999 11996
rect 20055 11994 20079 11996
rect 20135 11994 20141 11996
rect 19895 11942 19897 11994
rect 20077 11942 20079 11994
rect 19833 11940 19839 11942
rect 19895 11940 19919 11942
rect 19975 11940 19999 11942
rect 20055 11940 20079 11942
rect 20135 11940 20141 11942
rect 19833 11931 20141 11940
rect 27607 11996 27915 12005
rect 27607 11994 27613 11996
rect 27669 11994 27693 11996
rect 27749 11994 27773 11996
rect 27829 11994 27853 11996
rect 27909 11994 27915 11996
rect 27669 11942 27671 11994
rect 27851 11942 27853 11994
rect 27607 11940 27613 11942
rect 27669 11940 27693 11942
rect 27749 11940 27773 11942
rect 27829 11940 27853 11942
rect 27909 11940 27915 11942
rect 27607 11931 27915 11940
rect 8172 11452 8480 11461
rect 8172 11450 8178 11452
rect 8234 11450 8258 11452
rect 8314 11450 8338 11452
rect 8394 11450 8418 11452
rect 8474 11450 8480 11452
rect 8234 11398 8236 11450
rect 8416 11398 8418 11450
rect 8172 11396 8178 11398
rect 8234 11396 8258 11398
rect 8314 11396 8338 11398
rect 8394 11396 8418 11398
rect 8474 11396 8480 11398
rect 8172 11387 8480 11396
rect 15946 11452 16254 11461
rect 15946 11450 15952 11452
rect 16008 11450 16032 11452
rect 16088 11450 16112 11452
rect 16168 11450 16192 11452
rect 16248 11450 16254 11452
rect 16008 11398 16010 11450
rect 16190 11398 16192 11450
rect 15946 11396 15952 11398
rect 16008 11396 16032 11398
rect 16088 11396 16112 11398
rect 16168 11396 16192 11398
rect 16248 11396 16254 11398
rect 15946 11387 16254 11396
rect 23720 11452 24028 11461
rect 23720 11450 23726 11452
rect 23782 11450 23806 11452
rect 23862 11450 23886 11452
rect 23942 11450 23966 11452
rect 24022 11450 24028 11452
rect 23782 11398 23784 11450
rect 23964 11398 23966 11450
rect 23720 11396 23726 11398
rect 23782 11396 23806 11398
rect 23862 11396 23886 11398
rect 23942 11396 23966 11398
rect 24022 11396 24028 11398
rect 23720 11387 24028 11396
rect 31494 11452 31802 11461
rect 31494 11450 31500 11452
rect 31556 11450 31580 11452
rect 31636 11450 31660 11452
rect 31716 11450 31740 11452
rect 31796 11450 31802 11452
rect 31556 11398 31558 11450
rect 31738 11398 31740 11450
rect 31494 11396 31500 11398
rect 31556 11396 31580 11398
rect 31636 11396 31660 11398
rect 31716 11396 31740 11398
rect 31796 11396 31802 11398
rect 31494 11387 31802 11396
rect 4285 10908 4593 10917
rect 4285 10906 4291 10908
rect 4347 10906 4371 10908
rect 4427 10906 4451 10908
rect 4507 10906 4531 10908
rect 4587 10906 4593 10908
rect 4347 10854 4349 10906
rect 4529 10854 4531 10906
rect 4285 10852 4291 10854
rect 4347 10852 4371 10854
rect 4427 10852 4451 10854
rect 4507 10852 4531 10854
rect 4587 10852 4593 10854
rect 4285 10843 4593 10852
rect 12059 10908 12367 10917
rect 12059 10906 12065 10908
rect 12121 10906 12145 10908
rect 12201 10906 12225 10908
rect 12281 10906 12305 10908
rect 12361 10906 12367 10908
rect 12121 10854 12123 10906
rect 12303 10854 12305 10906
rect 12059 10852 12065 10854
rect 12121 10852 12145 10854
rect 12201 10852 12225 10854
rect 12281 10852 12305 10854
rect 12361 10852 12367 10854
rect 12059 10843 12367 10852
rect 19833 10908 20141 10917
rect 19833 10906 19839 10908
rect 19895 10906 19919 10908
rect 19975 10906 19999 10908
rect 20055 10906 20079 10908
rect 20135 10906 20141 10908
rect 19895 10854 19897 10906
rect 20077 10854 20079 10906
rect 19833 10852 19839 10854
rect 19895 10852 19919 10854
rect 19975 10852 19999 10854
rect 20055 10852 20079 10854
rect 20135 10852 20141 10854
rect 19833 10843 20141 10852
rect 27607 10908 27915 10917
rect 27607 10906 27613 10908
rect 27669 10906 27693 10908
rect 27749 10906 27773 10908
rect 27829 10906 27853 10908
rect 27909 10906 27915 10908
rect 27669 10854 27671 10906
rect 27851 10854 27853 10906
rect 27607 10852 27613 10854
rect 27669 10852 27693 10854
rect 27749 10852 27773 10854
rect 27829 10852 27853 10854
rect 27909 10852 27915 10854
rect 27607 10843 27915 10852
rect 8172 10364 8480 10373
rect 8172 10362 8178 10364
rect 8234 10362 8258 10364
rect 8314 10362 8338 10364
rect 8394 10362 8418 10364
rect 8474 10362 8480 10364
rect 8234 10310 8236 10362
rect 8416 10310 8418 10362
rect 8172 10308 8178 10310
rect 8234 10308 8258 10310
rect 8314 10308 8338 10310
rect 8394 10308 8418 10310
rect 8474 10308 8480 10310
rect 8172 10299 8480 10308
rect 15946 10364 16254 10373
rect 15946 10362 15952 10364
rect 16008 10362 16032 10364
rect 16088 10362 16112 10364
rect 16168 10362 16192 10364
rect 16248 10362 16254 10364
rect 16008 10310 16010 10362
rect 16190 10310 16192 10362
rect 15946 10308 15952 10310
rect 16008 10308 16032 10310
rect 16088 10308 16112 10310
rect 16168 10308 16192 10310
rect 16248 10308 16254 10310
rect 15946 10299 16254 10308
rect 23720 10364 24028 10373
rect 23720 10362 23726 10364
rect 23782 10362 23806 10364
rect 23862 10362 23886 10364
rect 23942 10362 23966 10364
rect 24022 10362 24028 10364
rect 23782 10310 23784 10362
rect 23964 10310 23966 10362
rect 23720 10308 23726 10310
rect 23782 10308 23806 10310
rect 23862 10308 23886 10310
rect 23942 10308 23966 10310
rect 24022 10308 24028 10310
rect 23720 10299 24028 10308
rect 31494 10364 31802 10373
rect 31494 10362 31500 10364
rect 31556 10362 31580 10364
rect 31636 10362 31660 10364
rect 31716 10362 31740 10364
rect 31796 10362 31802 10364
rect 31556 10310 31558 10362
rect 31738 10310 31740 10362
rect 31494 10308 31500 10310
rect 31556 10308 31580 10310
rect 31636 10308 31660 10310
rect 31716 10308 31740 10310
rect 31796 10308 31802 10310
rect 31494 10299 31802 10308
rect 4285 9820 4593 9829
rect 4285 9818 4291 9820
rect 4347 9818 4371 9820
rect 4427 9818 4451 9820
rect 4507 9818 4531 9820
rect 4587 9818 4593 9820
rect 4347 9766 4349 9818
rect 4529 9766 4531 9818
rect 4285 9764 4291 9766
rect 4347 9764 4371 9766
rect 4427 9764 4451 9766
rect 4507 9764 4531 9766
rect 4587 9764 4593 9766
rect 4285 9755 4593 9764
rect 12059 9820 12367 9829
rect 12059 9818 12065 9820
rect 12121 9818 12145 9820
rect 12201 9818 12225 9820
rect 12281 9818 12305 9820
rect 12361 9818 12367 9820
rect 12121 9766 12123 9818
rect 12303 9766 12305 9818
rect 12059 9764 12065 9766
rect 12121 9764 12145 9766
rect 12201 9764 12225 9766
rect 12281 9764 12305 9766
rect 12361 9764 12367 9766
rect 12059 9755 12367 9764
rect 19833 9820 20141 9829
rect 19833 9818 19839 9820
rect 19895 9818 19919 9820
rect 19975 9818 19999 9820
rect 20055 9818 20079 9820
rect 20135 9818 20141 9820
rect 19895 9766 19897 9818
rect 20077 9766 20079 9818
rect 19833 9764 19839 9766
rect 19895 9764 19919 9766
rect 19975 9764 19999 9766
rect 20055 9764 20079 9766
rect 20135 9764 20141 9766
rect 19833 9755 20141 9764
rect 27607 9820 27915 9829
rect 27607 9818 27613 9820
rect 27669 9818 27693 9820
rect 27749 9818 27773 9820
rect 27829 9818 27853 9820
rect 27909 9818 27915 9820
rect 27669 9766 27671 9818
rect 27851 9766 27853 9818
rect 27607 9764 27613 9766
rect 27669 9764 27693 9766
rect 27749 9764 27773 9766
rect 27829 9764 27853 9766
rect 27909 9764 27915 9766
rect 27607 9755 27915 9764
rect 8172 9276 8480 9285
rect 8172 9274 8178 9276
rect 8234 9274 8258 9276
rect 8314 9274 8338 9276
rect 8394 9274 8418 9276
rect 8474 9274 8480 9276
rect 8234 9222 8236 9274
rect 8416 9222 8418 9274
rect 8172 9220 8178 9222
rect 8234 9220 8258 9222
rect 8314 9220 8338 9222
rect 8394 9220 8418 9222
rect 8474 9220 8480 9222
rect 8172 9211 8480 9220
rect 15946 9276 16254 9285
rect 15946 9274 15952 9276
rect 16008 9274 16032 9276
rect 16088 9274 16112 9276
rect 16168 9274 16192 9276
rect 16248 9274 16254 9276
rect 16008 9222 16010 9274
rect 16190 9222 16192 9274
rect 15946 9220 15952 9222
rect 16008 9220 16032 9222
rect 16088 9220 16112 9222
rect 16168 9220 16192 9222
rect 16248 9220 16254 9222
rect 15946 9211 16254 9220
rect 23720 9276 24028 9285
rect 23720 9274 23726 9276
rect 23782 9274 23806 9276
rect 23862 9274 23886 9276
rect 23942 9274 23966 9276
rect 24022 9274 24028 9276
rect 23782 9222 23784 9274
rect 23964 9222 23966 9274
rect 23720 9220 23726 9222
rect 23782 9220 23806 9222
rect 23862 9220 23886 9222
rect 23942 9220 23966 9222
rect 24022 9220 24028 9222
rect 23720 9211 24028 9220
rect 31494 9276 31802 9285
rect 31494 9274 31500 9276
rect 31556 9274 31580 9276
rect 31636 9274 31660 9276
rect 31716 9274 31740 9276
rect 31796 9274 31802 9276
rect 31556 9222 31558 9274
rect 31738 9222 31740 9274
rect 31494 9220 31500 9222
rect 31556 9220 31580 9222
rect 31636 9220 31660 9222
rect 31716 9220 31740 9222
rect 31796 9220 31802 9222
rect 31494 9211 31802 9220
rect 4285 8732 4593 8741
rect 4285 8730 4291 8732
rect 4347 8730 4371 8732
rect 4427 8730 4451 8732
rect 4507 8730 4531 8732
rect 4587 8730 4593 8732
rect 4347 8678 4349 8730
rect 4529 8678 4531 8730
rect 4285 8676 4291 8678
rect 4347 8676 4371 8678
rect 4427 8676 4451 8678
rect 4507 8676 4531 8678
rect 4587 8676 4593 8678
rect 4285 8667 4593 8676
rect 12059 8732 12367 8741
rect 12059 8730 12065 8732
rect 12121 8730 12145 8732
rect 12201 8730 12225 8732
rect 12281 8730 12305 8732
rect 12361 8730 12367 8732
rect 12121 8678 12123 8730
rect 12303 8678 12305 8730
rect 12059 8676 12065 8678
rect 12121 8676 12145 8678
rect 12201 8676 12225 8678
rect 12281 8676 12305 8678
rect 12361 8676 12367 8678
rect 12059 8667 12367 8676
rect 19833 8732 20141 8741
rect 19833 8730 19839 8732
rect 19895 8730 19919 8732
rect 19975 8730 19999 8732
rect 20055 8730 20079 8732
rect 20135 8730 20141 8732
rect 19895 8678 19897 8730
rect 20077 8678 20079 8730
rect 19833 8676 19839 8678
rect 19895 8676 19919 8678
rect 19975 8676 19999 8678
rect 20055 8676 20079 8678
rect 20135 8676 20141 8678
rect 19833 8667 20141 8676
rect 27607 8732 27915 8741
rect 27607 8730 27613 8732
rect 27669 8730 27693 8732
rect 27749 8730 27773 8732
rect 27829 8730 27853 8732
rect 27909 8730 27915 8732
rect 27669 8678 27671 8730
rect 27851 8678 27853 8730
rect 27607 8676 27613 8678
rect 27669 8676 27693 8678
rect 27749 8676 27773 8678
rect 27829 8676 27853 8678
rect 27909 8676 27915 8678
rect 27607 8667 27915 8676
rect 8172 8188 8480 8197
rect 8172 8186 8178 8188
rect 8234 8186 8258 8188
rect 8314 8186 8338 8188
rect 8394 8186 8418 8188
rect 8474 8186 8480 8188
rect 8234 8134 8236 8186
rect 8416 8134 8418 8186
rect 8172 8132 8178 8134
rect 8234 8132 8258 8134
rect 8314 8132 8338 8134
rect 8394 8132 8418 8134
rect 8474 8132 8480 8134
rect 8172 8123 8480 8132
rect 15946 8188 16254 8197
rect 15946 8186 15952 8188
rect 16008 8186 16032 8188
rect 16088 8186 16112 8188
rect 16168 8186 16192 8188
rect 16248 8186 16254 8188
rect 16008 8134 16010 8186
rect 16190 8134 16192 8186
rect 15946 8132 15952 8134
rect 16008 8132 16032 8134
rect 16088 8132 16112 8134
rect 16168 8132 16192 8134
rect 16248 8132 16254 8134
rect 15946 8123 16254 8132
rect 23720 8188 24028 8197
rect 23720 8186 23726 8188
rect 23782 8186 23806 8188
rect 23862 8186 23886 8188
rect 23942 8186 23966 8188
rect 24022 8186 24028 8188
rect 23782 8134 23784 8186
rect 23964 8134 23966 8186
rect 23720 8132 23726 8134
rect 23782 8132 23806 8134
rect 23862 8132 23886 8134
rect 23942 8132 23966 8134
rect 24022 8132 24028 8134
rect 23720 8123 24028 8132
rect 31494 8188 31802 8197
rect 31494 8186 31500 8188
rect 31556 8186 31580 8188
rect 31636 8186 31660 8188
rect 31716 8186 31740 8188
rect 31796 8186 31802 8188
rect 31556 8134 31558 8186
rect 31738 8134 31740 8186
rect 31494 8132 31500 8134
rect 31556 8132 31580 8134
rect 31636 8132 31660 8134
rect 31716 8132 31740 8134
rect 31796 8132 31802 8134
rect 31494 8123 31802 8132
rect 4285 7644 4593 7653
rect 4285 7642 4291 7644
rect 4347 7642 4371 7644
rect 4427 7642 4451 7644
rect 4507 7642 4531 7644
rect 4587 7642 4593 7644
rect 4347 7590 4349 7642
rect 4529 7590 4531 7642
rect 4285 7588 4291 7590
rect 4347 7588 4371 7590
rect 4427 7588 4451 7590
rect 4507 7588 4531 7590
rect 4587 7588 4593 7590
rect 4285 7579 4593 7588
rect 12059 7644 12367 7653
rect 12059 7642 12065 7644
rect 12121 7642 12145 7644
rect 12201 7642 12225 7644
rect 12281 7642 12305 7644
rect 12361 7642 12367 7644
rect 12121 7590 12123 7642
rect 12303 7590 12305 7642
rect 12059 7588 12065 7590
rect 12121 7588 12145 7590
rect 12201 7588 12225 7590
rect 12281 7588 12305 7590
rect 12361 7588 12367 7590
rect 12059 7579 12367 7588
rect 19833 7644 20141 7653
rect 19833 7642 19839 7644
rect 19895 7642 19919 7644
rect 19975 7642 19999 7644
rect 20055 7642 20079 7644
rect 20135 7642 20141 7644
rect 19895 7590 19897 7642
rect 20077 7590 20079 7642
rect 19833 7588 19839 7590
rect 19895 7588 19919 7590
rect 19975 7588 19999 7590
rect 20055 7588 20079 7590
rect 20135 7588 20141 7590
rect 19833 7579 20141 7588
rect 27607 7644 27915 7653
rect 27607 7642 27613 7644
rect 27669 7642 27693 7644
rect 27749 7642 27773 7644
rect 27829 7642 27853 7644
rect 27909 7642 27915 7644
rect 27669 7590 27671 7642
rect 27851 7590 27853 7642
rect 27607 7588 27613 7590
rect 27669 7588 27693 7590
rect 27749 7588 27773 7590
rect 27829 7588 27853 7590
rect 27909 7588 27915 7590
rect 27607 7579 27915 7588
rect 8172 7100 8480 7109
rect 8172 7098 8178 7100
rect 8234 7098 8258 7100
rect 8314 7098 8338 7100
rect 8394 7098 8418 7100
rect 8474 7098 8480 7100
rect 8234 7046 8236 7098
rect 8416 7046 8418 7098
rect 8172 7044 8178 7046
rect 8234 7044 8258 7046
rect 8314 7044 8338 7046
rect 8394 7044 8418 7046
rect 8474 7044 8480 7046
rect 8172 7035 8480 7044
rect 15946 7100 16254 7109
rect 15946 7098 15952 7100
rect 16008 7098 16032 7100
rect 16088 7098 16112 7100
rect 16168 7098 16192 7100
rect 16248 7098 16254 7100
rect 16008 7046 16010 7098
rect 16190 7046 16192 7098
rect 15946 7044 15952 7046
rect 16008 7044 16032 7046
rect 16088 7044 16112 7046
rect 16168 7044 16192 7046
rect 16248 7044 16254 7046
rect 15946 7035 16254 7044
rect 23720 7100 24028 7109
rect 23720 7098 23726 7100
rect 23782 7098 23806 7100
rect 23862 7098 23886 7100
rect 23942 7098 23966 7100
rect 24022 7098 24028 7100
rect 23782 7046 23784 7098
rect 23964 7046 23966 7098
rect 23720 7044 23726 7046
rect 23782 7044 23806 7046
rect 23862 7044 23886 7046
rect 23942 7044 23966 7046
rect 24022 7044 24028 7046
rect 23720 7035 24028 7044
rect 31494 7100 31802 7109
rect 31494 7098 31500 7100
rect 31556 7098 31580 7100
rect 31636 7098 31660 7100
rect 31716 7098 31740 7100
rect 31796 7098 31802 7100
rect 31556 7046 31558 7098
rect 31738 7046 31740 7098
rect 31494 7044 31500 7046
rect 31556 7044 31580 7046
rect 31636 7044 31660 7046
rect 31716 7044 31740 7046
rect 31796 7044 31802 7046
rect 31494 7035 31802 7044
rect 4285 6556 4593 6565
rect 4285 6554 4291 6556
rect 4347 6554 4371 6556
rect 4427 6554 4451 6556
rect 4507 6554 4531 6556
rect 4587 6554 4593 6556
rect 4347 6502 4349 6554
rect 4529 6502 4531 6554
rect 4285 6500 4291 6502
rect 4347 6500 4371 6502
rect 4427 6500 4451 6502
rect 4507 6500 4531 6502
rect 4587 6500 4593 6502
rect 4285 6491 4593 6500
rect 12059 6556 12367 6565
rect 12059 6554 12065 6556
rect 12121 6554 12145 6556
rect 12201 6554 12225 6556
rect 12281 6554 12305 6556
rect 12361 6554 12367 6556
rect 12121 6502 12123 6554
rect 12303 6502 12305 6554
rect 12059 6500 12065 6502
rect 12121 6500 12145 6502
rect 12201 6500 12225 6502
rect 12281 6500 12305 6502
rect 12361 6500 12367 6502
rect 12059 6491 12367 6500
rect 19833 6556 20141 6565
rect 19833 6554 19839 6556
rect 19895 6554 19919 6556
rect 19975 6554 19999 6556
rect 20055 6554 20079 6556
rect 20135 6554 20141 6556
rect 19895 6502 19897 6554
rect 20077 6502 20079 6554
rect 19833 6500 19839 6502
rect 19895 6500 19919 6502
rect 19975 6500 19999 6502
rect 20055 6500 20079 6502
rect 20135 6500 20141 6502
rect 19833 6491 20141 6500
rect 27607 6556 27915 6565
rect 27607 6554 27613 6556
rect 27669 6554 27693 6556
rect 27749 6554 27773 6556
rect 27829 6554 27853 6556
rect 27909 6554 27915 6556
rect 27669 6502 27671 6554
rect 27851 6502 27853 6554
rect 27607 6500 27613 6502
rect 27669 6500 27693 6502
rect 27749 6500 27773 6502
rect 27829 6500 27853 6502
rect 27909 6500 27915 6502
rect 27607 6491 27915 6500
rect 8172 6012 8480 6021
rect 8172 6010 8178 6012
rect 8234 6010 8258 6012
rect 8314 6010 8338 6012
rect 8394 6010 8418 6012
rect 8474 6010 8480 6012
rect 8234 5958 8236 6010
rect 8416 5958 8418 6010
rect 8172 5956 8178 5958
rect 8234 5956 8258 5958
rect 8314 5956 8338 5958
rect 8394 5956 8418 5958
rect 8474 5956 8480 5958
rect 8172 5947 8480 5956
rect 15946 6012 16254 6021
rect 15946 6010 15952 6012
rect 16008 6010 16032 6012
rect 16088 6010 16112 6012
rect 16168 6010 16192 6012
rect 16248 6010 16254 6012
rect 16008 5958 16010 6010
rect 16190 5958 16192 6010
rect 15946 5956 15952 5958
rect 16008 5956 16032 5958
rect 16088 5956 16112 5958
rect 16168 5956 16192 5958
rect 16248 5956 16254 5958
rect 15946 5947 16254 5956
rect 23720 6012 24028 6021
rect 23720 6010 23726 6012
rect 23782 6010 23806 6012
rect 23862 6010 23886 6012
rect 23942 6010 23966 6012
rect 24022 6010 24028 6012
rect 23782 5958 23784 6010
rect 23964 5958 23966 6010
rect 23720 5956 23726 5958
rect 23782 5956 23806 5958
rect 23862 5956 23886 5958
rect 23942 5956 23966 5958
rect 24022 5956 24028 5958
rect 23720 5947 24028 5956
rect 31494 6012 31802 6021
rect 31494 6010 31500 6012
rect 31556 6010 31580 6012
rect 31636 6010 31660 6012
rect 31716 6010 31740 6012
rect 31796 6010 31802 6012
rect 31556 5958 31558 6010
rect 31738 5958 31740 6010
rect 31494 5956 31500 5958
rect 31556 5956 31580 5958
rect 31636 5956 31660 5958
rect 31716 5956 31740 5958
rect 31796 5956 31802 5958
rect 31494 5947 31802 5956
rect 4285 5468 4593 5477
rect 4285 5466 4291 5468
rect 4347 5466 4371 5468
rect 4427 5466 4451 5468
rect 4507 5466 4531 5468
rect 4587 5466 4593 5468
rect 4347 5414 4349 5466
rect 4529 5414 4531 5466
rect 4285 5412 4291 5414
rect 4347 5412 4371 5414
rect 4427 5412 4451 5414
rect 4507 5412 4531 5414
rect 4587 5412 4593 5414
rect 4285 5403 4593 5412
rect 12059 5468 12367 5477
rect 12059 5466 12065 5468
rect 12121 5466 12145 5468
rect 12201 5466 12225 5468
rect 12281 5466 12305 5468
rect 12361 5466 12367 5468
rect 12121 5414 12123 5466
rect 12303 5414 12305 5466
rect 12059 5412 12065 5414
rect 12121 5412 12145 5414
rect 12201 5412 12225 5414
rect 12281 5412 12305 5414
rect 12361 5412 12367 5414
rect 12059 5403 12367 5412
rect 19833 5468 20141 5477
rect 19833 5466 19839 5468
rect 19895 5466 19919 5468
rect 19975 5466 19999 5468
rect 20055 5466 20079 5468
rect 20135 5466 20141 5468
rect 19895 5414 19897 5466
rect 20077 5414 20079 5466
rect 19833 5412 19839 5414
rect 19895 5412 19919 5414
rect 19975 5412 19999 5414
rect 20055 5412 20079 5414
rect 20135 5412 20141 5414
rect 19833 5403 20141 5412
rect 27607 5468 27915 5477
rect 27607 5466 27613 5468
rect 27669 5466 27693 5468
rect 27749 5466 27773 5468
rect 27829 5466 27853 5468
rect 27909 5466 27915 5468
rect 27669 5414 27671 5466
rect 27851 5414 27853 5466
rect 27607 5412 27613 5414
rect 27669 5412 27693 5414
rect 27749 5412 27773 5414
rect 27829 5412 27853 5414
rect 27909 5412 27915 5414
rect 27607 5403 27915 5412
rect 8172 4924 8480 4933
rect 8172 4922 8178 4924
rect 8234 4922 8258 4924
rect 8314 4922 8338 4924
rect 8394 4922 8418 4924
rect 8474 4922 8480 4924
rect 8234 4870 8236 4922
rect 8416 4870 8418 4922
rect 8172 4868 8178 4870
rect 8234 4868 8258 4870
rect 8314 4868 8338 4870
rect 8394 4868 8418 4870
rect 8474 4868 8480 4870
rect 8172 4859 8480 4868
rect 15946 4924 16254 4933
rect 15946 4922 15952 4924
rect 16008 4922 16032 4924
rect 16088 4922 16112 4924
rect 16168 4922 16192 4924
rect 16248 4922 16254 4924
rect 16008 4870 16010 4922
rect 16190 4870 16192 4922
rect 15946 4868 15952 4870
rect 16008 4868 16032 4870
rect 16088 4868 16112 4870
rect 16168 4868 16192 4870
rect 16248 4868 16254 4870
rect 15946 4859 16254 4868
rect 23720 4924 24028 4933
rect 23720 4922 23726 4924
rect 23782 4922 23806 4924
rect 23862 4922 23886 4924
rect 23942 4922 23966 4924
rect 24022 4922 24028 4924
rect 23782 4870 23784 4922
rect 23964 4870 23966 4922
rect 23720 4868 23726 4870
rect 23782 4868 23806 4870
rect 23862 4868 23886 4870
rect 23942 4868 23966 4870
rect 24022 4868 24028 4870
rect 23720 4859 24028 4868
rect 31494 4924 31802 4933
rect 31494 4922 31500 4924
rect 31556 4922 31580 4924
rect 31636 4922 31660 4924
rect 31716 4922 31740 4924
rect 31796 4922 31802 4924
rect 31556 4870 31558 4922
rect 31738 4870 31740 4922
rect 31494 4868 31500 4870
rect 31556 4868 31580 4870
rect 31636 4868 31660 4870
rect 31716 4868 31740 4870
rect 31796 4868 31802 4870
rect 31494 4859 31802 4868
rect 4285 4380 4593 4389
rect 4285 4378 4291 4380
rect 4347 4378 4371 4380
rect 4427 4378 4451 4380
rect 4507 4378 4531 4380
rect 4587 4378 4593 4380
rect 4347 4326 4349 4378
rect 4529 4326 4531 4378
rect 4285 4324 4291 4326
rect 4347 4324 4371 4326
rect 4427 4324 4451 4326
rect 4507 4324 4531 4326
rect 4587 4324 4593 4326
rect 4285 4315 4593 4324
rect 12059 4380 12367 4389
rect 12059 4378 12065 4380
rect 12121 4378 12145 4380
rect 12201 4378 12225 4380
rect 12281 4378 12305 4380
rect 12361 4378 12367 4380
rect 12121 4326 12123 4378
rect 12303 4326 12305 4378
rect 12059 4324 12065 4326
rect 12121 4324 12145 4326
rect 12201 4324 12225 4326
rect 12281 4324 12305 4326
rect 12361 4324 12367 4326
rect 12059 4315 12367 4324
rect 19833 4380 20141 4389
rect 19833 4378 19839 4380
rect 19895 4378 19919 4380
rect 19975 4378 19999 4380
rect 20055 4378 20079 4380
rect 20135 4378 20141 4380
rect 19895 4326 19897 4378
rect 20077 4326 20079 4378
rect 19833 4324 19839 4326
rect 19895 4324 19919 4326
rect 19975 4324 19999 4326
rect 20055 4324 20079 4326
rect 20135 4324 20141 4326
rect 19833 4315 20141 4324
rect 27607 4380 27915 4389
rect 27607 4378 27613 4380
rect 27669 4378 27693 4380
rect 27749 4378 27773 4380
rect 27829 4378 27853 4380
rect 27909 4378 27915 4380
rect 27669 4326 27671 4378
rect 27851 4326 27853 4378
rect 27607 4324 27613 4326
rect 27669 4324 27693 4326
rect 27749 4324 27773 4326
rect 27829 4324 27853 4326
rect 27909 4324 27915 4326
rect 27607 4315 27915 4324
rect 8172 3836 8480 3845
rect 8172 3834 8178 3836
rect 8234 3834 8258 3836
rect 8314 3834 8338 3836
rect 8394 3834 8418 3836
rect 8474 3834 8480 3836
rect 8234 3782 8236 3834
rect 8416 3782 8418 3834
rect 8172 3780 8178 3782
rect 8234 3780 8258 3782
rect 8314 3780 8338 3782
rect 8394 3780 8418 3782
rect 8474 3780 8480 3782
rect 8172 3771 8480 3780
rect 15946 3836 16254 3845
rect 15946 3834 15952 3836
rect 16008 3834 16032 3836
rect 16088 3834 16112 3836
rect 16168 3834 16192 3836
rect 16248 3834 16254 3836
rect 16008 3782 16010 3834
rect 16190 3782 16192 3834
rect 15946 3780 15952 3782
rect 16008 3780 16032 3782
rect 16088 3780 16112 3782
rect 16168 3780 16192 3782
rect 16248 3780 16254 3782
rect 15946 3771 16254 3780
rect 23720 3836 24028 3845
rect 23720 3834 23726 3836
rect 23782 3834 23806 3836
rect 23862 3834 23886 3836
rect 23942 3834 23966 3836
rect 24022 3834 24028 3836
rect 23782 3782 23784 3834
rect 23964 3782 23966 3834
rect 23720 3780 23726 3782
rect 23782 3780 23806 3782
rect 23862 3780 23886 3782
rect 23942 3780 23966 3782
rect 24022 3780 24028 3782
rect 23720 3771 24028 3780
rect 31494 3836 31802 3845
rect 31494 3834 31500 3836
rect 31556 3834 31580 3836
rect 31636 3834 31660 3836
rect 31716 3834 31740 3836
rect 31796 3834 31802 3836
rect 31556 3782 31558 3834
rect 31738 3782 31740 3834
rect 31494 3780 31500 3782
rect 31556 3780 31580 3782
rect 31636 3780 31660 3782
rect 31716 3780 31740 3782
rect 31796 3780 31802 3782
rect 31494 3771 31802 3780
rect 4285 3292 4593 3301
rect 4285 3290 4291 3292
rect 4347 3290 4371 3292
rect 4427 3290 4451 3292
rect 4507 3290 4531 3292
rect 4587 3290 4593 3292
rect 4347 3238 4349 3290
rect 4529 3238 4531 3290
rect 4285 3236 4291 3238
rect 4347 3236 4371 3238
rect 4427 3236 4451 3238
rect 4507 3236 4531 3238
rect 4587 3236 4593 3238
rect 4285 3227 4593 3236
rect 12059 3292 12367 3301
rect 12059 3290 12065 3292
rect 12121 3290 12145 3292
rect 12201 3290 12225 3292
rect 12281 3290 12305 3292
rect 12361 3290 12367 3292
rect 12121 3238 12123 3290
rect 12303 3238 12305 3290
rect 12059 3236 12065 3238
rect 12121 3236 12145 3238
rect 12201 3236 12225 3238
rect 12281 3236 12305 3238
rect 12361 3236 12367 3238
rect 12059 3227 12367 3236
rect 19833 3292 20141 3301
rect 19833 3290 19839 3292
rect 19895 3290 19919 3292
rect 19975 3290 19999 3292
rect 20055 3290 20079 3292
rect 20135 3290 20141 3292
rect 19895 3238 19897 3290
rect 20077 3238 20079 3290
rect 19833 3236 19839 3238
rect 19895 3236 19919 3238
rect 19975 3236 19999 3238
rect 20055 3236 20079 3238
rect 20135 3236 20141 3238
rect 19833 3227 20141 3236
rect 27607 3292 27915 3301
rect 27607 3290 27613 3292
rect 27669 3290 27693 3292
rect 27749 3290 27773 3292
rect 27829 3290 27853 3292
rect 27909 3290 27915 3292
rect 27669 3238 27671 3290
rect 27851 3238 27853 3290
rect 27607 3236 27613 3238
rect 27669 3236 27693 3238
rect 27749 3236 27773 3238
rect 27829 3236 27853 3238
rect 27909 3236 27915 3238
rect 27607 3227 27915 3236
rect 8172 2748 8480 2757
rect 8172 2746 8178 2748
rect 8234 2746 8258 2748
rect 8314 2746 8338 2748
rect 8394 2746 8418 2748
rect 8474 2746 8480 2748
rect 8234 2694 8236 2746
rect 8416 2694 8418 2746
rect 8172 2692 8178 2694
rect 8234 2692 8258 2694
rect 8314 2692 8338 2694
rect 8394 2692 8418 2694
rect 8474 2692 8480 2694
rect 8172 2683 8480 2692
rect 15946 2748 16254 2757
rect 15946 2746 15952 2748
rect 16008 2746 16032 2748
rect 16088 2746 16112 2748
rect 16168 2746 16192 2748
rect 16248 2746 16254 2748
rect 16008 2694 16010 2746
rect 16190 2694 16192 2746
rect 15946 2692 15952 2694
rect 16008 2692 16032 2694
rect 16088 2692 16112 2694
rect 16168 2692 16192 2694
rect 16248 2692 16254 2694
rect 15946 2683 16254 2692
rect 23720 2748 24028 2757
rect 23720 2746 23726 2748
rect 23782 2746 23806 2748
rect 23862 2746 23886 2748
rect 23942 2746 23966 2748
rect 24022 2746 24028 2748
rect 23782 2694 23784 2746
rect 23964 2694 23966 2746
rect 23720 2692 23726 2694
rect 23782 2692 23806 2694
rect 23862 2692 23886 2694
rect 23942 2692 23966 2694
rect 24022 2692 24028 2694
rect 23720 2683 24028 2692
rect 31494 2748 31802 2757
rect 31494 2746 31500 2748
rect 31556 2746 31580 2748
rect 31636 2746 31660 2748
rect 31716 2746 31740 2748
rect 31796 2746 31802 2748
rect 31556 2694 31558 2746
rect 31738 2694 31740 2746
rect 31494 2692 31500 2694
rect 31556 2692 31580 2694
rect 31636 2692 31660 2694
rect 31716 2692 31740 2694
rect 31796 2692 31802 2694
rect 31494 2683 31802 2692
rect 4285 2204 4593 2213
rect 4285 2202 4291 2204
rect 4347 2202 4371 2204
rect 4427 2202 4451 2204
rect 4507 2202 4531 2204
rect 4587 2202 4593 2204
rect 4347 2150 4349 2202
rect 4529 2150 4531 2202
rect 4285 2148 4291 2150
rect 4347 2148 4371 2150
rect 4427 2148 4451 2150
rect 4507 2148 4531 2150
rect 4587 2148 4593 2150
rect 4285 2139 4593 2148
rect 12059 2204 12367 2213
rect 12059 2202 12065 2204
rect 12121 2202 12145 2204
rect 12201 2202 12225 2204
rect 12281 2202 12305 2204
rect 12361 2202 12367 2204
rect 12121 2150 12123 2202
rect 12303 2150 12305 2202
rect 12059 2148 12065 2150
rect 12121 2148 12145 2150
rect 12201 2148 12225 2150
rect 12281 2148 12305 2150
rect 12361 2148 12367 2150
rect 12059 2139 12367 2148
rect 19833 2204 20141 2213
rect 19833 2202 19839 2204
rect 19895 2202 19919 2204
rect 19975 2202 19999 2204
rect 20055 2202 20079 2204
rect 20135 2202 20141 2204
rect 19895 2150 19897 2202
rect 20077 2150 20079 2202
rect 19833 2148 19839 2150
rect 19895 2148 19919 2150
rect 19975 2148 19999 2150
rect 20055 2148 20079 2150
rect 20135 2148 20141 2150
rect 19833 2139 20141 2148
rect 27607 2204 27915 2213
rect 27607 2202 27613 2204
rect 27669 2202 27693 2204
rect 27749 2202 27773 2204
rect 27829 2202 27853 2204
rect 27909 2202 27915 2204
rect 27669 2150 27671 2202
rect 27851 2150 27853 2202
rect 27607 2148 27613 2150
rect 27669 2148 27693 2150
rect 27749 2148 27773 2150
rect 27829 2148 27853 2150
rect 27909 2148 27915 2150
rect 27607 2139 27915 2148
rect 8172 1660 8480 1669
rect 8172 1658 8178 1660
rect 8234 1658 8258 1660
rect 8314 1658 8338 1660
rect 8394 1658 8418 1660
rect 8474 1658 8480 1660
rect 8234 1606 8236 1658
rect 8416 1606 8418 1658
rect 8172 1604 8178 1606
rect 8234 1604 8258 1606
rect 8314 1604 8338 1606
rect 8394 1604 8418 1606
rect 8474 1604 8480 1606
rect 8172 1595 8480 1604
rect 15946 1660 16254 1669
rect 15946 1658 15952 1660
rect 16008 1658 16032 1660
rect 16088 1658 16112 1660
rect 16168 1658 16192 1660
rect 16248 1658 16254 1660
rect 16008 1606 16010 1658
rect 16190 1606 16192 1658
rect 15946 1604 15952 1606
rect 16008 1604 16032 1606
rect 16088 1604 16112 1606
rect 16168 1604 16192 1606
rect 16248 1604 16254 1606
rect 15946 1595 16254 1604
rect 23720 1660 24028 1669
rect 23720 1658 23726 1660
rect 23782 1658 23806 1660
rect 23862 1658 23886 1660
rect 23942 1658 23966 1660
rect 24022 1658 24028 1660
rect 23782 1606 23784 1658
rect 23964 1606 23966 1658
rect 23720 1604 23726 1606
rect 23782 1604 23806 1606
rect 23862 1604 23886 1606
rect 23942 1604 23966 1606
rect 24022 1604 24028 1606
rect 23720 1595 24028 1604
rect 31494 1660 31802 1669
rect 31494 1658 31500 1660
rect 31556 1658 31580 1660
rect 31636 1658 31660 1660
rect 31716 1658 31740 1660
rect 31796 1658 31802 1660
rect 31556 1606 31558 1658
rect 31738 1606 31740 1658
rect 31494 1604 31500 1606
rect 31556 1604 31580 1606
rect 31636 1604 31660 1606
rect 31716 1604 31740 1606
rect 31796 1604 31802 1606
rect 31494 1595 31802 1604
rect 4285 1116 4593 1125
rect 4285 1114 4291 1116
rect 4347 1114 4371 1116
rect 4427 1114 4451 1116
rect 4507 1114 4531 1116
rect 4587 1114 4593 1116
rect 4347 1062 4349 1114
rect 4529 1062 4531 1114
rect 4285 1060 4291 1062
rect 4347 1060 4371 1062
rect 4427 1060 4451 1062
rect 4507 1060 4531 1062
rect 4587 1060 4593 1062
rect 4285 1051 4593 1060
rect 12059 1116 12367 1125
rect 12059 1114 12065 1116
rect 12121 1114 12145 1116
rect 12201 1114 12225 1116
rect 12281 1114 12305 1116
rect 12361 1114 12367 1116
rect 12121 1062 12123 1114
rect 12303 1062 12305 1114
rect 12059 1060 12065 1062
rect 12121 1060 12145 1062
rect 12201 1060 12225 1062
rect 12281 1060 12305 1062
rect 12361 1060 12367 1062
rect 12059 1051 12367 1060
rect 19833 1116 20141 1125
rect 19833 1114 19839 1116
rect 19895 1114 19919 1116
rect 19975 1114 19999 1116
rect 20055 1114 20079 1116
rect 20135 1114 20141 1116
rect 19895 1062 19897 1114
rect 20077 1062 20079 1114
rect 19833 1060 19839 1062
rect 19895 1060 19919 1062
rect 19975 1060 19999 1062
rect 20055 1060 20079 1062
rect 20135 1060 20141 1062
rect 19833 1051 20141 1060
rect 27607 1116 27915 1125
rect 27607 1114 27613 1116
rect 27669 1114 27693 1116
rect 27749 1114 27773 1116
rect 27829 1114 27853 1116
rect 27909 1114 27915 1116
rect 27669 1062 27671 1114
rect 27851 1062 27853 1114
rect 27607 1060 27613 1062
rect 27669 1060 27693 1062
rect 27749 1060 27773 1062
rect 27829 1060 27853 1062
rect 27909 1060 27915 1062
rect 27607 1051 27915 1060
rect 8172 572 8480 581
rect 8172 570 8178 572
rect 8234 570 8258 572
rect 8314 570 8338 572
rect 8394 570 8418 572
rect 8474 570 8480 572
rect 8234 518 8236 570
rect 8416 518 8418 570
rect 8172 516 8178 518
rect 8234 516 8258 518
rect 8314 516 8338 518
rect 8394 516 8418 518
rect 8474 516 8480 518
rect 8172 507 8480 516
rect 15946 572 16254 581
rect 15946 570 15952 572
rect 16008 570 16032 572
rect 16088 570 16112 572
rect 16168 570 16192 572
rect 16248 570 16254 572
rect 16008 518 16010 570
rect 16190 518 16192 570
rect 15946 516 15952 518
rect 16008 516 16032 518
rect 16088 516 16112 518
rect 16168 516 16192 518
rect 16248 516 16254 518
rect 15946 507 16254 516
rect 23720 572 24028 581
rect 23720 570 23726 572
rect 23782 570 23806 572
rect 23862 570 23886 572
rect 23942 570 23966 572
rect 24022 570 24028 572
rect 23782 518 23784 570
rect 23964 518 23966 570
rect 23720 516 23726 518
rect 23782 516 23806 518
rect 23862 516 23886 518
rect 23942 516 23966 518
rect 24022 516 24028 518
rect 23720 507 24028 516
rect 31494 572 31802 581
rect 31494 570 31500 572
rect 31556 570 31580 572
rect 31636 570 31660 572
rect 31716 570 31740 572
rect 31796 570 31802 572
rect 31556 518 31558 570
rect 31738 518 31740 570
rect 31494 516 31500 518
rect 31556 516 31580 518
rect 31636 516 31660 518
rect 31716 516 31740 518
rect 31796 516 31802 518
rect 31494 507 31802 516
<< via2 >>
rect 29182 22208 29238 22264
rect 4526 21936 4582 21992
rect 846 21800 902 21856
rect 1582 21800 1638 21856
rect 2318 21800 2374 21856
rect 3238 21800 3294 21856
rect 3790 21800 3846 21856
rect 4291 21786 4347 21788
rect 4371 21786 4427 21788
rect 4451 21786 4507 21788
rect 4531 21786 4587 21788
rect 4291 21734 4337 21786
rect 4337 21734 4347 21786
rect 4371 21734 4401 21786
rect 4401 21734 4413 21786
rect 4413 21734 4427 21786
rect 4451 21734 4465 21786
rect 4465 21734 4477 21786
rect 4477 21734 4507 21786
rect 4531 21734 4541 21786
rect 4541 21734 4587 21786
rect 4291 21732 4347 21734
rect 4371 21732 4427 21734
rect 4451 21732 4507 21734
rect 4531 21732 4587 21734
rect 8390 21936 8446 21992
rect 16302 21936 16358 21992
rect 5262 21800 5318 21856
rect 5998 21800 6054 21856
rect 6734 21800 6790 21856
rect 7470 21800 7526 21856
rect 8942 21800 8998 21856
rect 9678 21800 9734 21856
rect 10414 21800 10470 21856
rect 11150 21800 11206 21856
rect 11886 21800 11942 21856
rect 12622 21800 12678 21856
rect 13542 21800 13598 21856
rect 14094 21800 14150 21856
rect 14830 21800 14886 21856
rect 15566 21800 15622 21856
rect 12065 21786 12121 21788
rect 12145 21786 12201 21788
rect 12225 21786 12281 21788
rect 12305 21786 12361 21788
rect 12065 21734 12111 21786
rect 12111 21734 12121 21786
rect 12145 21734 12175 21786
rect 12175 21734 12187 21786
rect 12187 21734 12201 21786
rect 12225 21734 12239 21786
rect 12239 21734 12251 21786
rect 12251 21734 12281 21786
rect 12305 21734 12315 21786
rect 12315 21734 12361 21786
rect 12065 21732 12121 21734
rect 12145 21732 12201 21734
rect 12225 21732 12281 21734
rect 12305 21732 12361 21734
rect 17038 21800 17094 21856
rect 19839 21786 19895 21788
rect 19919 21786 19975 21788
rect 19999 21786 20055 21788
rect 20079 21786 20135 21788
rect 19839 21734 19885 21786
rect 19885 21734 19895 21786
rect 19919 21734 19949 21786
rect 19949 21734 19961 21786
rect 19961 21734 19975 21786
rect 19999 21734 20013 21786
rect 20013 21734 20025 21786
rect 20025 21734 20055 21786
rect 20079 21734 20089 21786
rect 20089 21734 20135 21786
rect 19839 21732 19895 21734
rect 19919 21732 19975 21734
rect 19999 21732 20055 21734
rect 20079 21732 20135 21734
rect 27613 21786 27669 21788
rect 27693 21786 27749 21788
rect 27773 21786 27829 21788
rect 27853 21786 27909 21788
rect 27613 21734 27659 21786
rect 27659 21734 27669 21786
rect 27693 21734 27723 21786
rect 27723 21734 27735 21786
rect 27735 21734 27749 21786
rect 27773 21734 27787 21786
rect 27787 21734 27799 21786
rect 27799 21734 27829 21786
rect 27853 21734 27863 21786
rect 27863 21734 27909 21786
rect 27613 21732 27669 21734
rect 27693 21732 27749 21734
rect 27773 21732 27829 21734
rect 27853 21732 27909 21734
rect 29734 21800 29790 21856
rect 8178 21242 8234 21244
rect 8258 21242 8314 21244
rect 8338 21242 8394 21244
rect 8418 21242 8474 21244
rect 8178 21190 8224 21242
rect 8224 21190 8234 21242
rect 8258 21190 8288 21242
rect 8288 21190 8300 21242
rect 8300 21190 8314 21242
rect 8338 21190 8352 21242
rect 8352 21190 8364 21242
rect 8364 21190 8394 21242
rect 8418 21190 8428 21242
rect 8428 21190 8474 21242
rect 8178 21188 8234 21190
rect 8258 21188 8314 21190
rect 8338 21188 8394 21190
rect 8418 21188 8474 21190
rect 15952 21242 16008 21244
rect 16032 21242 16088 21244
rect 16112 21242 16168 21244
rect 16192 21242 16248 21244
rect 15952 21190 15998 21242
rect 15998 21190 16008 21242
rect 16032 21190 16062 21242
rect 16062 21190 16074 21242
rect 16074 21190 16088 21242
rect 16112 21190 16126 21242
rect 16126 21190 16138 21242
rect 16138 21190 16168 21242
rect 16192 21190 16202 21242
rect 16202 21190 16248 21242
rect 15952 21188 16008 21190
rect 16032 21188 16088 21190
rect 16112 21188 16168 21190
rect 16192 21188 16248 21190
rect 23726 21242 23782 21244
rect 23806 21242 23862 21244
rect 23886 21242 23942 21244
rect 23966 21242 24022 21244
rect 23726 21190 23772 21242
rect 23772 21190 23782 21242
rect 23806 21190 23836 21242
rect 23836 21190 23848 21242
rect 23848 21190 23862 21242
rect 23886 21190 23900 21242
rect 23900 21190 23912 21242
rect 23912 21190 23942 21242
rect 23966 21190 23976 21242
rect 23976 21190 24022 21242
rect 23726 21188 23782 21190
rect 23806 21188 23862 21190
rect 23886 21188 23942 21190
rect 23966 21188 24022 21190
rect 4291 20698 4347 20700
rect 4371 20698 4427 20700
rect 4451 20698 4507 20700
rect 4531 20698 4587 20700
rect 4291 20646 4337 20698
rect 4337 20646 4347 20698
rect 4371 20646 4401 20698
rect 4401 20646 4413 20698
rect 4413 20646 4427 20698
rect 4451 20646 4465 20698
rect 4465 20646 4477 20698
rect 4477 20646 4507 20698
rect 4531 20646 4541 20698
rect 4541 20646 4587 20698
rect 4291 20644 4347 20646
rect 4371 20644 4427 20646
rect 4451 20644 4507 20646
rect 4531 20644 4587 20646
rect 12065 20698 12121 20700
rect 12145 20698 12201 20700
rect 12225 20698 12281 20700
rect 12305 20698 12361 20700
rect 12065 20646 12111 20698
rect 12111 20646 12121 20698
rect 12145 20646 12175 20698
rect 12175 20646 12187 20698
rect 12187 20646 12201 20698
rect 12225 20646 12239 20698
rect 12239 20646 12251 20698
rect 12251 20646 12281 20698
rect 12305 20646 12315 20698
rect 12315 20646 12361 20698
rect 12065 20644 12121 20646
rect 12145 20644 12201 20646
rect 12225 20644 12281 20646
rect 12305 20644 12361 20646
rect 19839 20698 19895 20700
rect 19919 20698 19975 20700
rect 19999 20698 20055 20700
rect 20079 20698 20135 20700
rect 19839 20646 19885 20698
rect 19885 20646 19895 20698
rect 19919 20646 19949 20698
rect 19949 20646 19961 20698
rect 19961 20646 19975 20698
rect 19999 20646 20013 20698
rect 20013 20646 20025 20698
rect 20025 20646 20055 20698
rect 20079 20646 20089 20698
rect 20089 20646 20135 20698
rect 19839 20644 19895 20646
rect 19919 20644 19975 20646
rect 19999 20644 20055 20646
rect 20079 20644 20135 20646
rect 8178 20154 8234 20156
rect 8258 20154 8314 20156
rect 8338 20154 8394 20156
rect 8418 20154 8474 20156
rect 8178 20102 8224 20154
rect 8224 20102 8234 20154
rect 8258 20102 8288 20154
rect 8288 20102 8300 20154
rect 8300 20102 8314 20154
rect 8338 20102 8352 20154
rect 8352 20102 8364 20154
rect 8364 20102 8394 20154
rect 8418 20102 8428 20154
rect 8428 20102 8474 20154
rect 8178 20100 8234 20102
rect 8258 20100 8314 20102
rect 8338 20100 8394 20102
rect 8418 20100 8474 20102
rect 15952 20154 16008 20156
rect 16032 20154 16088 20156
rect 16112 20154 16168 20156
rect 16192 20154 16248 20156
rect 15952 20102 15998 20154
rect 15998 20102 16008 20154
rect 16032 20102 16062 20154
rect 16062 20102 16074 20154
rect 16074 20102 16088 20154
rect 16112 20102 16126 20154
rect 16126 20102 16138 20154
rect 16138 20102 16168 20154
rect 16192 20102 16202 20154
rect 16202 20102 16248 20154
rect 15952 20100 16008 20102
rect 16032 20100 16088 20102
rect 16112 20100 16168 20102
rect 16192 20100 16248 20102
rect 23726 20154 23782 20156
rect 23806 20154 23862 20156
rect 23886 20154 23942 20156
rect 23966 20154 24022 20156
rect 23726 20102 23772 20154
rect 23772 20102 23782 20154
rect 23806 20102 23836 20154
rect 23836 20102 23848 20154
rect 23848 20102 23862 20154
rect 23886 20102 23900 20154
rect 23900 20102 23912 20154
rect 23912 20102 23942 20154
rect 23966 20102 23976 20154
rect 23976 20102 24022 20154
rect 23726 20100 23782 20102
rect 23806 20100 23862 20102
rect 23886 20100 23942 20102
rect 23966 20100 24022 20102
rect 4291 19610 4347 19612
rect 4371 19610 4427 19612
rect 4451 19610 4507 19612
rect 4531 19610 4587 19612
rect 4291 19558 4337 19610
rect 4337 19558 4347 19610
rect 4371 19558 4401 19610
rect 4401 19558 4413 19610
rect 4413 19558 4427 19610
rect 4451 19558 4465 19610
rect 4465 19558 4477 19610
rect 4477 19558 4507 19610
rect 4531 19558 4541 19610
rect 4541 19558 4587 19610
rect 4291 19556 4347 19558
rect 4371 19556 4427 19558
rect 4451 19556 4507 19558
rect 4531 19556 4587 19558
rect 12065 19610 12121 19612
rect 12145 19610 12201 19612
rect 12225 19610 12281 19612
rect 12305 19610 12361 19612
rect 12065 19558 12111 19610
rect 12111 19558 12121 19610
rect 12145 19558 12175 19610
rect 12175 19558 12187 19610
rect 12187 19558 12201 19610
rect 12225 19558 12239 19610
rect 12239 19558 12251 19610
rect 12251 19558 12281 19610
rect 12305 19558 12315 19610
rect 12315 19558 12361 19610
rect 12065 19556 12121 19558
rect 12145 19556 12201 19558
rect 12225 19556 12281 19558
rect 12305 19556 12361 19558
rect 19839 19610 19895 19612
rect 19919 19610 19975 19612
rect 19999 19610 20055 19612
rect 20079 19610 20135 19612
rect 19839 19558 19885 19610
rect 19885 19558 19895 19610
rect 19919 19558 19949 19610
rect 19949 19558 19961 19610
rect 19961 19558 19975 19610
rect 19999 19558 20013 19610
rect 20013 19558 20025 19610
rect 20025 19558 20055 19610
rect 20079 19558 20089 19610
rect 20089 19558 20135 19610
rect 19839 19556 19895 19558
rect 19919 19556 19975 19558
rect 19999 19556 20055 19558
rect 20079 19556 20135 19558
rect 31500 21242 31556 21244
rect 31580 21242 31636 21244
rect 31660 21242 31716 21244
rect 31740 21242 31796 21244
rect 31500 21190 31546 21242
rect 31546 21190 31556 21242
rect 31580 21190 31610 21242
rect 31610 21190 31622 21242
rect 31622 21190 31636 21242
rect 31660 21190 31674 21242
rect 31674 21190 31686 21242
rect 31686 21190 31716 21242
rect 31740 21190 31750 21242
rect 31750 21190 31796 21242
rect 31500 21188 31556 21190
rect 31580 21188 31636 21190
rect 31660 21188 31716 21190
rect 31740 21188 31796 21190
rect 27613 20698 27669 20700
rect 27693 20698 27749 20700
rect 27773 20698 27829 20700
rect 27853 20698 27909 20700
rect 27613 20646 27659 20698
rect 27659 20646 27669 20698
rect 27693 20646 27723 20698
rect 27723 20646 27735 20698
rect 27735 20646 27749 20698
rect 27773 20646 27787 20698
rect 27787 20646 27799 20698
rect 27799 20646 27829 20698
rect 27853 20646 27863 20698
rect 27863 20646 27909 20698
rect 27613 20644 27669 20646
rect 27693 20644 27749 20646
rect 27773 20644 27829 20646
rect 27853 20644 27909 20646
rect 31500 20154 31556 20156
rect 31580 20154 31636 20156
rect 31660 20154 31716 20156
rect 31740 20154 31796 20156
rect 31500 20102 31546 20154
rect 31546 20102 31556 20154
rect 31580 20102 31610 20154
rect 31610 20102 31622 20154
rect 31622 20102 31636 20154
rect 31660 20102 31674 20154
rect 31674 20102 31686 20154
rect 31686 20102 31716 20154
rect 31740 20102 31750 20154
rect 31750 20102 31796 20154
rect 31500 20100 31556 20102
rect 31580 20100 31636 20102
rect 31660 20100 31716 20102
rect 31740 20100 31796 20102
rect 27613 19610 27669 19612
rect 27693 19610 27749 19612
rect 27773 19610 27829 19612
rect 27853 19610 27909 19612
rect 27613 19558 27659 19610
rect 27659 19558 27669 19610
rect 27693 19558 27723 19610
rect 27723 19558 27735 19610
rect 27735 19558 27749 19610
rect 27773 19558 27787 19610
rect 27787 19558 27799 19610
rect 27799 19558 27829 19610
rect 27853 19558 27863 19610
rect 27863 19558 27909 19610
rect 27613 19556 27669 19558
rect 27693 19556 27749 19558
rect 27773 19556 27829 19558
rect 27853 19556 27909 19558
rect 25686 19216 25742 19272
rect 8178 19066 8234 19068
rect 8258 19066 8314 19068
rect 8338 19066 8394 19068
rect 8418 19066 8474 19068
rect 8178 19014 8224 19066
rect 8224 19014 8234 19066
rect 8258 19014 8288 19066
rect 8288 19014 8300 19066
rect 8300 19014 8314 19066
rect 8338 19014 8352 19066
rect 8352 19014 8364 19066
rect 8364 19014 8394 19066
rect 8418 19014 8428 19066
rect 8428 19014 8474 19066
rect 8178 19012 8234 19014
rect 8258 19012 8314 19014
rect 8338 19012 8394 19014
rect 8418 19012 8474 19014
rect 15952 19066 16008 19068
rect 16032 19066 16088 19068
rect 16112 19066 16168 19068
rect 16192 19066 16248 19068
rect 15952 19014 15998 19066
rect 15998 19014 16008 19066
rect 16032 19014 16062 19066
rect 16062 19014 16074 19066
rect 16074 19014 16088 19066
rect 16112 19014 16126 19066
rect 16126 19014 16138 19066
rect 16138 19014 16168 19066
rect 16192 19014 16202 19066
rect 16202 19014 16248 19066
rect 15952 19012 16008 19014
rect 16032 19012 16088 19014
rect 16112 19012 16168 19014
rect 16192 19012 16248 19014
rect 23726 19066 23782 19068
rect 23806 19066 23862 19068
rect 23886 19066 23942 19068
rect 23966 19066 24022 19068
rect 23726 19014 23772 19066
rect 23772 19014 23782 19066
rect 23806 19014 23836 19066
rect 23836 19014 23848 19066
rect 23848 19014 23862 19066
rect 23886 19014 23900 19066
rect 23900 19014 23912 19066
rect 23912 19014 23942 19066
rect 23966 19014 23976 19066
rect 23976 19014 24022 19066
rect 23726 19012 23782 19014
rect 23806 19012 23862 19014
rect 23886 19012 23942 19014
rect 23966 19012 24022 19014
rect 31500 19066 31556 19068
rect 31580 19066 31636 19068
rect 31660 19066 31716 19068
rect 31740 19066 31796 19068
rect 31500 19014 31546 19066
rect 31546 19014 31556 19066
rect 31580 19014 31610 19066
rect 31610 19014 31622 19066
rect 31622 19014 31636 19066
rect 31660 19014 31674 19066
rect 31674 19014 31686 19066
rect 31686 19014 31716 19066
rect 31740 19014 31750 19066
rect 31750 19014 31796 19066
rect 31500 19012 31556 19014
rect 31580 19012 31636 19014
rect 31660 19012 31716 19014
rect 31740 19012 31796 19014
rect 4291 18522 4347 18524
rect 4371 18522 4427 18524
rect 4451 18522 4507 18524
rect 4531 18522 4587 18524
rect 4291 18470 4337 18522
rect 4337 18470 4347 18522
rect 4371 18470 4401 18522
rect 4401 18470 4413 18522
rect 4413 18470 4427 18522
rect 4451 18470 4465 18522
rect 4465 18470 4477 18522
rect 4477 18470 4507 18522
rect 4531 18470 4541 18522
rect 4541 18470 4587 18522
rect 4291 18468 4347 18470
rect 4371 18468 4427 18470
rect 4451 18468 4507 18470
rect 4531 18468 4587 18470
rect 12065 18522 12121 18524
rect 12145 18522 12201 18524
rect 12225 18522 12281 18524
rect 12305 18522 12361 18524
rect 12065 18470 12111 18522
rect 12111 18470 12121 18522
rect 12145 18470 12175 18522
rect 12175 18470 12187 18522
rect 12187 18470 12201 18522
rect 12225 18470 12239 18522
rect 12239 18470 12251 18522
rect 12251 18470 12281 18522
rect 12305 18470 12315 18522
rect 12315 18470 12361 18522
rect 12065 18468 12121 18470
rect 12145 18468 12201 18470
rect 12225 18468 12281 18470
rect 12305 18468 12361 18470
rect 19839 18522 19895 18524
rect 19919 18522 19975 18524
rect 19999 18522 20055 18524
rect 20079 18522 20135 18524
rect 19839 18470 19885 18522
rect 19885 18470 19895 18522
rect 19919 18470 19949 18522
rect 19949 18470 19961 18522
rect 19961 18470 19975 18522
rect 19999 18470 20013 18522
rect 20013 18470 20025 18522
rect 20025 18470 20055 18522
rect 20079 18470 20089 18522
rect 20089 18470 20135 18522
rect 19839 18468 19895 18470
rect 19919 18468 19975 18470
rect 19999 18468 20055 18470
rect 20079 18468 20135 18470
rect 27613 18522 27669 18524
rect 27693 18522 27749 18524
rect 27773 18522 27829 18524
rect 27853 18522 27909 18524
rect 27613 18470 27659 18522
rect 27659 18470 27669 18522
rect 27693 18470 27723 18522
rect 27723 18470 27735 18522
rect 27735 18470 27749 18522
rect 27773 18470 27787 18522
rect 27787 18470 27799 18522
rect 27799 18470 27829 18522
rect 27853 18470 27863 18522
rect 27863 18470 27909 18522
rect 27613 18468 27669 18470
rect 27693 18468 27749 18470
rect 27773 18468 27829 18470
rect 27853 18468 27909 18470
rect 8178 17978 8234 17980
rect 8258 17978 8314 17980
rect 8338 17978 8394 17980
rect 8418 17978 8474 17980
rect 8178 17926 8224 17978
rect 8224 17926 8234 17978
rect 8258 17926 8288 17978
rect 8288 17926 8300 17978
rect 8300 17926 8314 17978
rect 8338 17926 8352 17978
rect 8352 17926 8364 17978
rect 8364 17926 8394 17978
rect 8418 17926 8428 17978
rect 8428 17926 8474 17978
rect 8178 17924 8234 17926
rect 8258 17924 8314 17926
rect 8338 17924 8394 17926
rect 8418 17924 8474 17926
rect 15952 17978 16008 17980
rect 16032 17978 16088 17980
rect 16112 17978 16168 17980
rect 16192 17978 16248 17980
rect 15952 17926 15998 17978
rect 15998 17926 16008 17978
rect 16032 17926 16062 17978
rect 16062 17926 16074 17978
rect 16074 17926 16088 17978
rect 16112 17926 16126 17978
rect 16126 17926 16138 17978
rect 16138 17926 16168 17978
rect 16192 17926 16202 17978
rect 16202 17926 16248 17978
rect 15952 17924 16008 17926
rect 16032 17924 16088 17926
rect 16112 17924 16168 17926
rect 16192 17924 16248 17926
rect 23726 17978 23782 17980
rect 23806 17978 23862 17980
rect 23886 17978 23942 17980
rect 23966 17978 24022 17980
rect 23726 17926 23772 17978
rect 23772 17926 23782 17978
rect 23806 17926 23836 17978
rect 23836 17926 23848 17978
rect 23848 17926 23862 17978
rect 23886 17926 23900 17978
rect 23900 17926 23912 17978
rect 23912 17926 23942 17978
rect 23966 17926 23976 17978
rect 23976 17926 24022 17978
rect 23726 17924 23782 17926
rect 23806 17924 23862 17926
rect 23886 17924 23942 17926
rect 23966 17924 24022 17926
rect 31500 17978 31556 17980
rect 31580 17978 31636 17980
rect 31660 17978 31716 17980
rect 31740 17978 31796 17980
rect 31500 17926 31546 17978
rect 31546 17926 31556 17978
rect 31580 17926 31610 17978
rect 31610 17926 31622 17978
rect 31622 17926 31636 17978
rect 31660 17926 31674 17978
rect 31674 17926 31686 17978
rect 31686 17926 31716 17978
rect 31740 17926 31750 17978
rect 31750 17926 31796 17978
rect 31500 17924 31556 17926
rect 31580 17924 31636 17926
rect 31660 17924 31716 17926
rect 31740 17924 31796 17926
rect 4291 17434 4347 17436
rect 4371 17434 4427 17436
rect 4451 17434 4507 17436
rect 4531 17434 4587 17436
rect 4291 17382 4337 17434
rect 4337 17382 4347 17434
rect 4371 17382 4401 17434
rect 4401 17382 4413 17434
rect 4413 17382 4427 17434
rect 4451 17382 4465 17434
rect 4465 17382 4477 17434
rect 4477 17382 4507 17434
rect 4531 17382 4541 17434
rect 4541 17382 4587 17434
rect 4291 17380 4347 17382
rect 4371 17380 4427 17382
rect 4451 17380 4507 17382
rect 4531 17380 4587 17382
rect 12065 17434 12121 17436
rect 12145 17434 12201 17436
rect 12225 17434 12281 17436
rect 12305 17434 12361 17436
rect 12065 17382 12111 17434
rect 12111 17382 12121 17434
rect 12145 17382 12175 17434
rect 12175 17382 12187 17434
rect 12187 17382 12201 17434
rect 12225 17382 12239 17434
rect 12239 17382 12251 17434
rect 12251 17382 12281 17434
rect 12305 17382 12315 17434
rect 12315 17382 12361 17434
rect 12065 17380 12121 17382
rect 12145 17380 12201 17382
rect 12225 17380 12281 17382
rect 12305 17380 12361 17382
rect 19839 17434 19895 17436
rect 19919 17434 19975 17436
rect 19999 17434 20055 17436
rect 20079 17434 20135 17436
rect 19839 17382 19885 17434
rect 19885 17382 19895 17434
rect 19919 17382 19949 17434
rect 19949 17382 19961 17434
rect 19961 17382 19975 17434
rect 19999 17382 20013 17434
rect 20013 17382 20025 17434
rect 20025 17382 20055 17434
rect 20079 17382 20089 17434
rect 20089 17382 20135 17434
rect 19839 17380 19895 17382
rect 19919 17380 19975 17382
rect 19999 17380 20055 17382
rect 20079 17380 20135 17382
rect 27613 17434 27669 17436
rect 27693 17434 27749 17436
rect 27773 17434 27829 17436
rect 27853 17434 27909 17436
rect 27613 17382 27659 17434
rect 27659 17382 27669 17434
rect 27693 17382 27723 17434
rect 27723 17382 27735 17434
rect 27735 17382 27749 17434
rect 27773 17382 27787 17434
rect 27787 17382 27799 17434
rect 27799 17382 27829 17434
rect 27853 17382 27863 17434
rect 27863 17382 27909 17434
rect 27613 17380 27669 17382
rect 27693 17380 27749 17382
rect 27773 17380 27829 17382
rect 27853 17380 27909 17382
rect 8178 16890 8234 16892
rect 8258 16890 8314 16892
rect 8338 16890 8394 16892
rect 8418 16890 8474 16892
rect 8178 16838 8224 16890
rect 8224 16838 8234 16890
rect 8258 16838 8288 16890
rect 8288 16838 8300 16890
rect 8300 16838 8314 16890
rect 8338 16838 8352 16890
rect 8352 16838 8364 16890
rect 8364 16838 8394 16890
rect 8418 16838 8428 16890
rect 8428 16838 8474 16890
rect 8178 16836 8234 16838
rect 8258 16836 8314 16838
rect 8338 16836 8394 16838
rect 8418 16836 8474 16838
rect 15952 16890 16008 16892
rect 16032 16890 16088 16892
rect 16112 16890 16168 16892
rect 16192 16890 16248 16892
rect 15952 16838 15998 16890
rect 15998 16838 16008 16890
rect 16032 16838 16062 16890
rect 16062 16838 16074 16890
rect 16074 16838 16088 16890
rect 16112 16838 16126 16890
rect 16126 16838 16138 16890
rect 16138 16838 16168 16890
rect 16192 16838 16202 16890
rect 16202 16838 16248 16890
rect 15952 16836 16008 16838
rect 16032 16836 16088 16838
rect 16112 16836 16168 16838
rect 16192 16836 16248 16838
rect 23726 16890 23782 16892
rect 23806 16890 23862 16892
rect 23886 16890 23942 16892
rect 23966 16890 24022 16892
rect 23726 16838 23772 16890
rect 23772 16838 23782 16890
rect 23806 16838 23836 16890
rect 23836 16838 23848 16890
rect 23848 16838 23862 16890
rect 23886 16838 23900 16890
rect 23900 16838 23912 16890
rect 23912 16838 23942 16890
rect 23966 16838 23976 16890
rect 23976 16838 24022 16890
rect 23726 16836 23782 16838
rect 23806 16836 23862 16838
rect 23886 16836 23942 16838
rect 23966 16836 24022 16838
rect 31500 16890 31556 16892
rect 31580 16890 31636 16892
rect 31660 16890 31716 16892
rect 31740 16890 31796 16892
rect 31500 16838 31546 16890
rect 31546 16838 31556 16890
rect 31580 16838 31610 16890
rect 31610 16838 31622 16890
rect 31622 16838 31636 16890
rect 31660 16838 31674 16890
rect 31674 16838 31686 16890
rect 31686 16838 31716 16890
rect 31740 16838 31750 16890
rect 31750 16838 31796 16890
rect 31500 16836 31556 16838
rect 31580 16836 31636 16838
rect 31660 16836 31716 16838
rect 31740 16836 31796 16838
rect 4291 16346 4347 16348
rect 4371 16346 4427 16348
rect 4451 16346 4507 16348
rect 4531 16346 4587 16348
rect 4291 16294 4337 16346
rect 4337 16294 4347 16346
rect 4371 16294 4401 16346
rect 4401 16294 4413 16346
rect 4413 16294 4427 16346
rect 4451 16294 4465 16346
rect 4465 16294 4477 16346
rect 4477 16294 4507 16346
rect 4531 16294 4541 16346
rect 4541 16294 4587 16346
rect 4291 16292 4347 16294
rect 4371 16292 4427 16294
rect 4451 16292 4507 16294
rect 4531 16292 4587 16294
rect 12065 16346 12121 16348
rect 12145 16346 12201 16348
rect 12225 16346 12281 16348
rect 12305 16346 12361 16348
rect 12065 16294 12111 16346
rect 12111 16294 12121 16346
rect 12145 16294 12175 16346
rect 12175 16294 12187 16346
rect 12187 16294 12201 16346
rect 12225 16294 12239 16346
rect 12239 16294 12251 16346
rect 12251 16294 12281 16346
rect 12305 16294 12315 16346
rect 12315 16294 12361 16346
rect 12065 16292 12121 16294
rect 12145 16292 12201 16294
rect 12225 16292 12281 16294
rect 12305 16292 12361 16294
rect 19839 16346 19895 16348
rect 19919 16346 19975 16348
rect 19999 16346 20055 16348
rect 20079 16346 20135 16348
rect 19839 16294 19885 16346
rect 19885 16294 19895 16346
rect 19919 16294 19949 16346
rect 19949 16294 19961 16346
rect 19961 16294 19975 16346
rect 19999 16294 20013 16346
rect 20013 16294 20025 16346
rect 20025 16294 20055 16346
rect 20079 16294 20089 16346
rect 20089 16294 20135 16346
rect 19839 16292 19895 16294
rect 19919 16292 19975 16294
rect 19999 16292 20055 16294
rect 20079 16292 20135 16294
rect 27613 16346 27669 16348
rect 27693 16346 27749 16348
rect 27773 16346 27829 16348
rect 27853 16346 27909 16348
rect 27613 16294 27659 16346
rect 27659 16294 27669 16346
rect 27693 16294 27723 16346
rect 27723 16294 27735 16346
rect 27735 16294 27749 16346
rect 27773 16294 27787 16346
rect 27787 16294 27799 16346
rect 27799 16294 27829 16346
rect 27853 16294 27863 16346
rect 27863 16294 27909 16346
rect 27613 16292 27669 16294
rect 27693 16292 27749 16294
rect 27773 16292 27829 16294
rect 27853 16292 27909 16294
rect 8178 15802 8234 15804
rect 8258 15802 8314 15804
rect 8338 15802 8394 15804
rect 8418 15802 8474 15804
rect 8178 15750 8224 15802
rect 8224 15750 8234 15802
rect 8258 15750 8288 15802
rect 8288 15750 8300 15802
rect 8300 15750 8314 15802
rect 8338 15750 8352 15802
rect 8352 15750 8364 15802
rect 8364 15750 8394 15802
rect 8418 15750 8428 15802
rect 8428 15750 8474 15802
rect 8178 15748 8234 15750
rect 8258 15748 8314 15750
rect 8338 15748 8394 15750
rect 8418 15748 8474 15750
rect 15952 15802 16008 15804
rect 16032 15802 16088 15804
rect 16112 15802 16168 15804
rect 16192 15802 16248 15804
rect 15952 15750 15998 15802
rect 15998 15750 16008 15802
rect 16032 15750 16062 15802
rect 16062 15750 16074 15802
rect 16074 15750 16088 15802
rect 16112 15750 16126 15802
rect 16126 15750 16138 15802
rect 16138 15750 16168 15802
rect 16192 15750 16202 15802
rect 16202 15750 16248 15802
rect 15952 15748 16008 15750
rect 16032 15748 16088 15750
rect 16112 15748 16168 15750
rect 16192 15748 16248 15750
rect 23726 15802 23782 15804
rect 23806 15802 23862 15804
rect 23886 15802 23942 15804
rect 23966 15802 24022 15804
rect 23726 15750 23772 15802
rect 23772 15750 23782 15802
rect 23806 15750 23836 15802
rect 23836 15750 23848 15802
rect 23848 15750 23862 15802
rect 23886 15750 23900 15802
rect 23900 15750 23912 15802
rect 23912 15750 23942 15802
rect 23966 15750 23976 15802
rect 23976 15750 24022 15802
rect 23726 15748 23782 15750
rect 23806 15748 23862 15750
rect 23886 15748 23942 15750
rect 23966 15748 24022 15750
rect 31500 15802 31556 15804
rect 31580 15802 31636 15804
rect 31660 15802 31716 15804
rect 31740 15802 31796 15804
rect 31500 15750 31546 15802
rect 31546 15750 31556 15802
rect 31580 15750 31610 15802
rect 31610 15750 31622 15802
rect 31622 15750 31636 15802
rect 31660 15750 31674 15802
rect 31674 15750 31686 15802
rect 31686 15750 31716 15802
rect 31740 15750 31750 15802
rect 31750 15750 31796 15802
rect 31500 15748 31556 15750
rect 31580 15748 31636 15750
rect 31660 15748 31716 15750
rect 31740 15748 31796 15750
rect 4291 15258 4347 15260
rect 4371 15258 4427 15260
rect 4451 15258 4507 15260
rect 4531 15258 4587 15260
rect 4291 15206 4337 15258
rect 4337 15206 4347 15258
rect 4371 15206 4401 15258
rect 4401 15206 4413 15258
rect 4413 15206 4427 15258
rect 4451 15206 4465 15258
rect 4465 15206 4477 15258
rect 4477 15206 4507 15258
rect 4531 15206 4541 15258
rect 4541 15206 4587 15258
rect 4291 15204 4347 15206
rect 4371 15204 4427 15206
rect 4451 15204 4507 15206
rect 4531 15204 4587 15206
rect 12065 15258 12121 15260
rect 12145 15258 12201 15260
rect 12225 15258 12281 15260
rect 12305 15258 12361 15260
rect 12065 15206 12111 15258
rect 12111 15206 12121 15258
rect 12145 15206 12175 15258
rect 12175 15206 12187 15258
rect 12187 15206 12201 15258
rect 12225 15206 12239 15258
rect 12239 15206 12251 15258
rect 12251 15206 12281 15258
rect 12305 15206 12315 15258
rect 12315 15206 12361 15258
rect 12065 15204 12121 15206
rect 12145 15204 12201 15206
rect 12225 15204 12281 15206
rect 12305 15204 12361 15206
rect 19839 15258 19895 15260
rect 19919 15258 19975 15260
rect 19999 15258 20055 15260
rect 20079 15258 20135 15260
rect 19839 15206 19885 15258
rect 19885 15206 19895 15258
rect 19919 15206 19949 15258
rect 19949 15206 19961 15258
rect 19961 15206 19975 15258
rect 19999 15206 20013 15258
rect 20013 15206 20025 15258
rect 20025 15206 20055 15258
rect 20079 15206 20089 15258
rect 20089 15206 20135 15258
rect 19839 15204 19895 15206
rect 19919 15204 19975 15206
rect 19999 15204 20055 15206
rect 20079 15204 20135 15206
rect 27613 15258 27669 15260
rect 27693 15258 27749 15260
rect 27773 15258 27829 15260
rect 27853 15258 27909 15260
rect 27613 15206 27659 15258
rect 27659 15206 27669 15258
rect 27693 15206 27723 15258
rect 27723 15206 27735 15258
rect 27735 15206 27749 15258
rect 27773 15206 27787 15258
rect 27787 15206 27799 15258
rect 27799 15206 27829 15258
rect 27853 15206 27863 15258
rect 27863 15206 27909 15258
rect 27613 15204 27669 15206
rect 27693 15204 27749 15206
rect 27773 15204 27829 15206
rect 27853 15204 27909 15206
rect 8178 14714 8234 14716
rect 8258 14714 8314 14716
rect 8338 14714 8394 14716
rect 8418 14714 8474 14716
rect 8178 14662 8224 14714
rect 8224 14662 8234 14714
rect 8258 14662 8288 14714
rect 8288 14662 8300 14714
rect 8300 14662 8314 14714
rect 8338 14662 8352 14714
rect 8352 14662 8364 14714
rect 8364 14662 8394 14714
rect 8418 14662 8428 14714
rect 8428 14662 8474 14714
rect 8178 14660 8234 14662
rect 8258 14660 8314 14662
rect 8338 14660 8394 14662
rect 8418 14660 8474 14662
rect 15952 14714 16008 14716
rect 16032 14714 16088 14716
rect 16112 14714 16168 14716
rect 16192 14714 16248 14716
rect 15952 14662 15998 14714
rect 15998 14662 16008 14714
rect 16032 14662 16062 14714
rect 16062 14662 16074 14714
rect 16074 14662 16088 14714
rect 16112 14662 16126 14714
rect 16126 14662 16138 14714
rect 16138 14662 16168 14714
rect 16192 14662 16202 14714
rect 16202 14662 16248 14714
rect 15952 14660 16008 14662
rect 16032 14660 16088 14662
rect 16112 14660 16168 14662
rect 16192 14660 16248 14662
rect 23726 14714 23782 14716
rect 23806 14714 23862 14716
rect 23886 14714 23942 14716
rect 23966 14714 24022 14716
rect 23726 14662 23772 14714
rect 23772 14662 23782 14714
rect 23806 14662 23836 14714
rect 23836 14662 23848 14714
rect 23848 14662 23862 14714
rect 23886 14662 23900 14714
rect 23900 14662 23912 14714
rect 23912 14662 23942 14714
rect 23966 14662 23976 14714
rect 23976 14662 24022 14714
rect 23726 14660 23782 14662
rect 23806 14660 23862 14662
rect 23886 14660 23942 14662
rect 23966 14660 24022 14662
rect 31500 14714 31556 14716
rect 31580 14714 31636 14716
rect 31660 14714 31716 14716
rect 31740 14714 31796 14716
rect 31500 14662 31546 14714
rect 31546 14662 31556 14714
rect 31580 14662 31610 14714
rect 31610 14662 31622 14714
rect 31622 14662 31636 14714
rect 31660 14662 31674 14714
rect 31674 14662 31686 14714
rect 31686 14662 31716 14714
rect 31740 14662 31750 14714
rect 31750 14662 31796 14714
rect 31500 14660 31556 14662
rect 31580 14660 31636 14662
rect 31660 14660 31716 14662
rect 31740 14660 31796 14662
rect 4291 14170 4347 14172
rect 4371 14170 4427 14172
rect 4451 14170 4507 14172
rect 4531 14170 4587 14172
rect 4291 14118 4337 14170
rect 4337 14118 4347 14170
rect 4371 14118 4401 14170
rect 4401 14118 4413 14170
rect 4413 14118 4427 14170
rect 4451 14118 4465 14170
rect 4465 14118 4477 14170
rect 4477 14118 4507 14170
rect 4531 14118 4541 14170
rect 4541 14118 4587 14170
rect 4291 14116 4347 14118
rect 4371 14116 4427 14118
rect 4451 14116 4507 14118
rect 4531 14116 4587 14118
rect 12065 14170 12121 14172
rect 12145 14170 12201 14172
rect 12225 14170 12281 14172
rect 12305 14170 12361 14172
rect 12065 14118 12111 14170
rect 12111 14118 12121 14170
rect 12145 14118 12175 14170
rect 12175 14118 12187 14170
rect 12187 14118 12201 14170
rect 12225 14118 12239 14170
rect 12239 14118 12251 14170
rect 12251 14118 12281 14170
rect 12305 14118 12315 14170
rect 12315 14118 12361 14170
rect 12065 14116 12121 14118
rect 12145 14116 12201 14118
rect 12225 14116 12281 14118
rect 12305 14116 12361 14118
rect 19839 14170 19895 14172
rect 19919 14170 19975 14172
rect 19999 14170 20055 14172
rect 20079 14170 20135 14172
rect 19839 14118 19885 14170
rect 19885 14118 19895 14170
rect 19919 14118 19949 14170
rect 19949 14118 19961 14170
rect 19961 14118 19975 14170
rect 19999 14118 20013 14170
rect 20013 14118 20025 14170
rect 20025 14118 20055 14170
rect 20079 14118 20089 14170
rect 20089 14118 20135 14170
rect 19839 14116 19895 14118
rect 19919 14116 19975 14118
rect 19999 14116 20055 14118
rect 20079 14116 20135 14118
rect 27613 14170 27669 14172
rect 27693 14170 27749 14172
rect 27773 14170 27829 14172
rect 27853 14170 27909 14172
rect 27613 14118 27659 14170
rect 27659 14118 27669 14170
rect 27693 14118 27723 14170
rect 27723 14118 27735 14170
rect 27735 14118 27749 14170
rect 27773 14118 27787 14170
rect 27787 14118 27799 14170
rect 27799 14118 27829 14170
rect 27853 14118 27863 14170
rect 27863 14118 27909 14170
rect 27613 14116 27669 14118
rect 27693 14116 27749 14118
rect 27773 14116 27829 14118
rect 27853 14116 27909 14118
rect 8178 13626 8234 13628
rect 8258 13626 8314 13628
rect 8338 13626 8394 13628
rect 8418 13626 8474 13628
rect 8178 13574 8224 13626
rect 8224 13574 8234 13626
rect 8258 13574 8288 13626
rect 8288 13574 8300 13626
rect 8300 13574 8314 13626
rect 8338 13574 8352 13626
rect 8352 13574 8364 13626
rect 8364 13574 8394 13626
rect 8418 13574 8428 13626
rect 8428 13574 8474 13626
rect 8178 13572 8234 13574
rect 8258 13572 8314 13574
rect 8338 13572 8394 13574
rect 8418 13572 8474 13574
rect 15952 13626 16008 13628
rect 16032 13626 16088 13628
rect 16112 13626 16168 13628
rect 16192 13626 16248 13628
rect 15952 13574 15998 13626
rect 15998 13574 16008 13626
rect 16032 13574 16062 13626
rect 16062 13574 16074 13626
rect 16074 13574 16088 13626
rect 16112 13574 16126 13626
rect 16126 13574 16138 13626
rect 16138 13574 16168 13626
rect 16192 13574 16202 13626
rect 16202 13574 16248 13626
rect 15952 13572 16008 13574
rect 16032 13572 16088 13574
rect 16112 13572 16168 13574
rect 16192 13572 16248 13574
rect 23726 13626 23782 13628
rect 23806 13626 23862 13628
rect 23886 13626 23942 13628
rect 23966 13626 24022 13628
rect 23726 13574 23772 13626
rect 23772 13574 23782 13626
rect 23806 13574 23836 13626
rect 23836 13574 23848 13626
rect 23848 13574 23862 13626
rect 23886 13574 23900 13626
rect 23900 13574 23912 13626
rect 23912 13574 23942 13626
rect 23966 13574 23976 13626
rect 23976 13574 24022 13626
rect 23726 13572 23782 13574
rect 23806 13572 23862 13574
rect 23886 13572 23942 13574
rect 23966 13572 24022 13574
rect 31500 13626 31556 13628
rect 31580 13626 31636 13628
rect 31660 13626 31716 13628
rect 31740 13626 31796 13628
rect 31500 13574 31546 13626
rect 31546 13574 31556 13626
rect 31580 13574 31610 13626
rect 31610 13574 31622 13626
rect 31622 13574 31636 13626
rect 31660 13574 31674 13626
rect 31674 13574 31686 13626
rect 31686 13574 31716 13626
rect 31740 13574 31750 13626
rect 31750 13574 31796 13626
rect 31500 13572 31556 13574
rect 31580 13572 31636 13574
rect 31660 13572 31716 13574
rect 31740 13572 31796 13574
rect 4291 13082 4347 13084
rect 4371 13082 4427 13084
rect 4451 13082 4507 13084
rect 4531 13082 4587 13084
rect 4291 13030 4337 13082
rect 4337 13030 4347 13082
rect 4371 13030 4401 13082
rect 4401 13030 4413 13082
rect 4413 13030 4427 13082
rect 4451 13030 4465 13082
rect 4465 13030 4477 13082
rect 4477 13030 4507 13082
rect 4531 13030 4541 13082
rect 4541 13030 4587 13082
rect 4291 13028 4347 13030
rect 4371 13028 4427 13030
rect 4451 13028 4507 13030
rect 4531 13028 4587 13030
rect 12065 13082 12121 13084
rect 12145 13082 12201 13084
rect 12225 13082 12281 13084
rect 12305 13082 12361 13084
rect 12065 13030 12111 13082
rect 12111 13030 12121 13082
rect 12145 13030 12175 13082
rect 12175 13030 12187 13082
rect 12187 13030 12201 13082
rect 12225 13030 12239 13082
rect 12239 13030 12251 13082
rect 12251 13030 12281 13082
rect 12305 13030 12315 13082
rect 12315 13030 12361 13082
rect 12065 13028 12121 13030
rect 12145 13028 12201 13030
rect 12225 13028 12281 13030
rect 12305 13028 12361 13030
rect 19839 13082 19895 13084
rect 19919 13082 19975 13084
rect 19999 13082 20055 13084
rect 20079 13082 20135 13084
rect 19839 13030 19885 13082
rect 19885 13030 19895 13082
rect 19919 13030 19949 13082
rect 19949 13030 19961 13082
rect 19961 13030 19975 13082
rect 19999 13030 20013 13082
rect 20013 13030 20025 13082
rect 20025 13030 20055 13082
rect 20079 13030 20089 13082
rect 20089 13030 20135 13082
rect 19839 13028 19895 13030
rect 19919 13028 19975 13030
rect 19999 13028 20055 13030
rect 20079 13028 20135 13030
rect 27613 13082 27669 13084
rect 27693 13082 27749 13084
rect 27773 13082 27829 13084
rect 27853 13082 27909 13084
rect 27613 13030 27659 13082
rect 27659 13030 27669 13082
rect 27693 13030 27723 13082
rect 27723 13030 27735 13082
rect 27735 13030 27749 13082
rect 27773 13030 27787 13082
rect 27787 13030 27799 13082
rect 27799 13030 27829 13082
rect 27853 13030 27863 13082
rect 27863 13030 27909 13082
rect 27613 13028 27669 13030
rect 27693 13028 27749 13030
rect 27773 13028 27829 13030
rect 27853 13028 27909 13030
rect 8178 12538 8234 12540
rect 8258 12538 8314 12540
rect 8338 12538 8394 12540
rect 8418 12538 8474 12540
rect 8178 12486 8224 12538
rect 8224 12486 8234 12538
rect 8258 12486 8288 12538
rect 8288 12486 8300 12538
rect 8300 12486 8314 12538
rect 8338 12486 8352 12538
rect 8352 12486 8364 12538
rect 8364 12486 8394 12538
rect 8418 12486 8428 12538
rect 8428 12486 8474 12538
rect 8178 12484 8234 12486
rect 8258 12484 8314 12486
rect 8338 12484 8394 12486
rect 8418 12484 8474 12486
rect 15952 12538 16008 12540
rect 16032 12538 16088 12540
rect 16112 12538 16168 12540
rect 16192 12538 16248 12540
rect 15952 12486 15998 12538
rect 15998 12486 16008 12538
rect 16032 12486 16062 12538
rect 16062 12486 16074 12538
rect 16074 12486 16088 12538
rect 16112 12486 16126 12538
rect 16126 12486 16138 12538
rect 16138 12486 16168 12538
rect 16192 12486 16202 12538
rect 16202 12486 16248 12538
rect 15952 12484 16008 12486
rect 16032 12484 16088 12486
rect 16112 12484 16168 12486
rect 16192 12484 16248 12486
rect 23726 12538 23782 12540
rect 23806 12538 23862 12540
rect 23886 12538 23942 12540
rect 23966 12538 24022 12540
rect 23726 12486 23772 12538
rect 23772 12486 23782 12538
rect 23806 12486 23836 12538
rect 23836 12486 23848 12538
rect 23848 12486 23862 12538
rect 23886 12486 23900 12538
rect 23900 12486 23912 12538
rect 23912 12486 23942 12538
rect 23966 12486 23976 12538
rect 23976 12486 24022 12538
rect 23726 12484 23782 12486
rect 23806 12484 23862 12486
rect 23886 12484 23942 12486
rect 23966 12484 24022 12486
rect 31500 12538 31556 12540
rect 31580 12538 31636 12540
rect 31660 12538 31716 12540
rect 31740 12538 31796 12540
rect 31500 12486 31546 12538
rect 31546 12486 31556 12538
rect 31580 12486 31610 12538
rect 31610 12486 31622 12538
rect 31622 12486 31636 12538
rect 31660 12486 31674 12538
rect 31674 12486 31686 12538
rect 31686 12486 31716 12538
rect 31740 12486 31750 12538
rect 31750 12486 31796 12538
rect 31500 12484 31556 12486
rect 31580 12484 31636 12486
rect 31660 12484 31716 12486
rect 31740 12484 31796 12486
rect 4291 11994 4347 11996
rect 4371 11994 4427 11996
rect 4451 11994 4507 11996
rect 4531 11994 4587 11996
rect 4291 11942 4337 11994
rect 4337 11942 4347 11994
rect 4371 11942 4401 11994
rect 4401 11942 4413 11994
rect 4413 11942 4427 11994
rect 4451 11942 4465 11994
rect 4465 11942 4477 11994
rect 4477 11942 4507 11994
rect 4531 11942 4541 11994
rect 4541 11942 4587 11994
rect 4291 11940 4347 11942
rect 4371 11940 4427 11942
rect 4451 11940 4507 11942
rect 4531 11940 4587 11942
rect 12065 11994 12121 11996
rect 12145 11994 12201 11996
rect 12225 11994 12281 11996
rect 12305 11994 12361 11996
rect 12065 11942 12111 11994
rect 12111 11942 12121 11994
rect 12145 11942 12175 11994
rect 12175 11942 12187 11994
rect 12187 11942 12201 11994
rect 12225 11942 12239 11994
rect 12239 11942 12251 11994
rect 12251 11942 12281 11994
rect 12305 11942 12315 11994
rect 12315 11942 12361 11994
rect 12065 11940 12121 11942
rect 12145 11940 12201 11942
rect 12225 11940 12281 11942
rect 12305 11940 12361 11942
rect 19839 11994 19895 11996
rect 19919 11994 19975 11996
rect 19999 11994 20055 11996
rect 20079 11994 20135 11996
rect 19839 11942 19885 11994
rect 19885 11942 19895 11994
rect 19919 11942 19949 11994
rect 19949 11942 19961 11994
rect 19961 11942 19975 11994
rect 19999 11942 20013 11994
rect 20013 11942 20025 11994
rect 20025 11942 20055 11994
rect 20079 11942 20089 11994
rect 20089 11942 20135 11994
rect 19839 11940 19895 11942
rect 19919 11940 19975 11942
rect 19999 11940 20055 11942
rect 20079 11940 20135 11942
rect 27613 11994 27669 11996
rect 27693 11994 27749 11996
rect 27773 11994 27829 11996
rect 27853 11994 27909 11996
rect 27613 11942 27659 11994
rect 27659 11942 27669 11994
rect 27693 11942 27723 11994
rect 27723 11942 27735 11994
rect 27735 11942 27749 11994
rect 27773 11942 27787 11994
rect 27787 11942 27799 11994
rect 27799 11942 27829 11994
rect 27853 11942 27863 11994
rect 27863 11942 27909 11994
rect 27613 11940 27669 11942
rect 27693 11940 27749 11942
rect 27773 11940 27829 11942
rect 27853 11940 27909 11942
rect 8178 11450 8234 11452
rect 8258 11450 8314 11452
rect 8338 11450 8394 11452
rect 8418 11450 8474 11452
rect 8178 11398 8224 11450
rect 8224 11398 8234 11450
rect 8258 11398 8288 11450
rect 8288 11398 8300 11450
rect 8300 11398 8314 11450
rect 8338 11398 8352 11450
rect 8352 11398 8364 11450
rect 8364 11398 8394 11450
rect 8418 11398 8428 11450
rect 8428 11398 8474 11450
rect 8178 11396 8234 11398
rect 8258 11396 8314 11398
rect 8338 11396 8394 11398
rect 8418 11396 8474 11398
rect 15952 11450 16008 11452
rect 16032 11450 16088 11452
rect 16112 11450 16168 11452
rect 16192 11450 16248 11452
rect 15952 11398 15998 11450
rect 15998 11398 16008 11450
rect 16032 11398 16062 11450
rect 16062 11398 16074 11450
rect 16074 11398 16088 11450
rect 16112 11398 16126 11450
rect 16126 11398 16138 11450
rect 16138 11398 16168 11450
rect 16192 11398 16202 11450
rect 16202 11398 16248 11450
rect 15952 11396 16008 11398
rect 16032 11396 16088 11398
rect 16112 11396 16168 11398
rect 16192 11396 16248 11398
rect 23726 11450 23782 11452
rect 23806 11450 23862 11452
rect 23886 11450 23942 11452
rect 23966 11450 24022 11452
rect 23726 11398 23772 11450
rect 23772 11398 23782 11450
rect 23806 11398 23836 11450
rect 23836 11398 23848 11450
rect 23848 11398 23862 11450
rect 23886 11398 23900 11450
rect 23900 11398 23912 11450
rect 23912 11398 23942 11450
rect 23966 11398 23976 11450
rect 23976 11398 24022 11450
rect 23726 11396 23782 11398
rect 23806 11396 23862 11398
rect 23886 11396 23942 11398
rect 23966 11396 24022 11398
rect 31500 11450 31556 11452
rect 31580 11450 31636 11452
rect 31660 11450 31716 11452
rect 31740 11450 31796 11452
rect 31500 11398 31546 11450
rect 31546 11398 31556 11450
rect 31580 11398 31610 11450
rect 31610 11398 31622 11450
rect 31622 11398 31636 11450
rect 31660 11398 31674 11450
rect 31674 11398 31686 11450
rect 31686 11398 31716 11450
rect 31740 11398 31750 11450
rect 31750 11398 31796 11450
rect 31500 11396 31556 11398
rect 31580 11396 31636 11398
rect 31660 11396 31716 11398
rect 31740 11396 31796 11398
rect 4291 10906 4347 10908
rect 4371 10906 4427 10908
rect 4451 10906 4507 10908
rect 4531 10906 4587 10908
rect 4291 10854 4337 10906
rect 4337 10854 4347 10906
rect 4371 10854 4401 10906
rect 4401 10854 4413 10906
rect 4413 10854 4427 10906
rect 4451 10854 4465 10906
rect 4465 10854 4477 10906
rect 4477 10854 4507 10906
rect 4531 10854 4541 10906
rect 4541 10854 4587 10906
rect 4291 10852 4347 10854
rect 4371 10852 4427 10854
rect 4451 10852 4507 10854
rect 4531 10852 4587 10854
rect 12065 10906 12121 10908
rect 12145 10906 12201 10908
rect 12225 10906 12281 10908
rect 12305 10906 12361 10908
rect 12065 10854 12111 10906
rect 12111 10854 12121 10906
rect 12145 10854 12175 10906
rect 12175 10854 12187 10906
rect 12187 10854 12201 10906
rect 12225 10854 12239 10906
rect 12239 10854 12251 10906
rect 12251 10854 12281 10906
rect 12305 10854 12315 10906
rect 12315 10854 12361 10906
rect 12065 10852 12121 10854
rect 12145 10852 12201 10854
rect 12225 10852 12281 10854
rect 12305 10852 12361 10854
rect 19839 10906 19895 10908
rect 19919 10906 19975 10908
rect 19999 10906 20055 10908
rect 20079 10906 20135 10908
rect 19839 10854 19885 10906
rect 19885 10854 19895 10906
rect 19919 10854 19949 10906
rect 19949 10854 19961 10906
rect 19961 10854 19975 10906
rect 19999 10854 20013 10906
rect 20013 10854 20025 10906
rect 20025 10854 20055 10906
rect 20079 10854 20089 10906
rect 20089 10854 20135 10906
rect 19839 10852 19895 10854
rect 19919 10852 19975 10854
rect 19999 10852 20055 10854
rect 20079 10852 20135 10854
rect 27613 10906 27669 10908
rect 27693 10906 27749 10908
rect 27773 10906 27829 10908
rect 27853 10906 27909 10908
rect 27613 10854 27659 10906
rect 27659 10854 27669 10906
rect 27693 10854 27723 10906
rect 27723 10854 27735 10906
rect 27735 10854 27749 10906
rect 27773 10854 27787 10906
rect 27787 10854 27799 10906
rect 27799 10854 27829 10906
rect 27853 10854 27863 10906
rect 27863 10854 27909 10906
rect 27613 10852 27669 10854
rect 27693 10852 27749 10854
rect 27773 10852 27829 10854
rect 27853 10852 27909 10854
rect 8178 10362 8234 10364
rect 8258 10362 8314 10364
rect 8338 10362 8394 10364
rect 8418 10362 8474 10364
rect 8178 10310 8224 10362
rect 8224 10310 8234 10362
rect 8258 10310 8288 10362
rect 8288 10310 8300 10362
rect 8300 10310 8314 10362
rect 8338 10310 8352 10362
rect 8352 10310 8364 10362
rect 8364 10310 8394 10362
rect 8418 10310 8428 10362
rect 8428 10310 8474 10362
rect 8178 10308 8234 10310
rect 8258 10308 8314 10310
rect 8338 10308 8394 10310
rect 8418 10308 8474 10310
rect 15952 10362 16008 10364
rect 16032 10362 16088 10364
rect 16112 10362 16168 10364
rect 16192 10362 16248 10364
rect 15952 10310 15998 10362
rect 15998 10310 16008 10362
rect 16032 10310 16062 10362
rect 16062 10310 16074 10362
rect 16074 10310 16088 10362
rect 16112 10310 16126 10362
rect 16126 10310 16138 10362
rect 16138 10310 16168 10362
rect 16192 10310 16202 10362
rect 16202 10310 16248 10362
rect 15952 10308 16008 10310
rect 16032 10308 16088 10310
rect 16112 10308 16168 10310
rect 16192 10308 16248 10310
rect 23726 10362 23782 10364
rect 23806 10362 23862 10364
rect 23886 10362 23942 10364
rect 23966 10362 24022 10364
rect 23726 10310 23772 10362
rect 23772 10310 23782 10362
rect 23806 10310 23836 10362
rect 23836 10310 23848 10362
rect 23848 10310 23862 10362
rect 23886 10310 23900 10362
rect 23900 10310 23912 10362
rect 23912 10310 23942 10362
rect 23966 10310 23976 10362
rect 23976 10310 24022 10362
rect 23726 10308 23782 10310
rect 23806 10308 23862 10310
rect 23886 10308 23942 10310
rect 23966 10308 24022 10310
rect 31500 10362 31556 10364
rect 31580 10362 31636 10364
rect 31660 10362 31716 10364
rect 31740 10362 31796 10364
rect 31500 10310 31546 10362
rect 31546 10310 31556 10362
rect 31580 10310 31610 10362
rect 31610 10310 31622 10362
rect 31622 10310 31636 10362
rect 31660 10310 31674 10362
rect 31674 10310 31686 10362
rect 31686 10310 31716 10362
rect 31740 10310 31750 10362
rect 31750 10310 31796 10362
rect 31500 10308 31556 10310
rect 31580 10308 31636 10310
rect 31660 10308 31716 10310
rect 31740 10308 31796 10310
rect 4291 9818 4347 9820
rect 4371 9818 4427 9820
rect 4451 9818 4507 9820
rect 4531 9818 4587 9820
rect 4291 9766 4337 9818
rect 4337 9766 4347 9818
rect 4371 9766 4401 9818
rect 4401 9766 4413 9818
rect 4413 9766 4427 9818
rect 4451 9766 4465 9818
rect 4465 9766 4477 9818
rect 4477 9766 4507 9818
rect 4531 9766 4541 9818
rect 4541 9766 4587 9818
rect 4291 9764 4347 9766
rect 4371 9764 4427 9766
rect 4451 9764 4507 9766
rect 4531 9764 4587 9766
rect 12065 9818 12121 9820
rect 12145 9818 12201 9820
rect 12225 9818 12281 9820
rect 12305 9818 12361 9820
rect 12065 9766 12111 9818
rect 12111 9766 12121 9818
rect 12145 9766 12175 9818
rect 12175 9766 12187 9818
rect 12187 9766 12201 9818
rect 12225 9766 12239 9818
rect 12239 9766 12251 9818
rect 12251 9766 12281 9818
rect 12305 9766 12315 9818
rect 12315 9766 12361 9818
rect 12065 9764 12121 9766
rect 12145 9764 12201 9766
rect 12225 9764 12281 9766
rect 12305 9764 12361 9766
rect 19839 9818 19895 9820
rect 19919 9818 19975 9820
rect 19999 9818 20055 9820
rect 20079 9818 20135 9820
rect 19839 9766 19885 9818
rect 19885 9766 19895 9818
rect 19919 9766 19949 9818
rect 19949 9766 19961 9818
rect 19961 9766 19975 9818
rect 19999 9766 20013 9818
rect 20013 9766 20025 9818
rect 20025 9766 20055 9818
rect 20079 9766 20089 9818
rect 20089 9766 20135 9818
rect 19839 9764 19895 9766
rect 19919 9764 19975 9766
rect 19999 9764 20055 9766
rect 20079 9764 20135 9766
rect 27613 9818 27669 9820
rect 27693 9818 27749 9820
rect 27773 9818 27829 9820
rect 27853 9818 27909 9820
rect 27613 9766 27659 9818
rect 27659 9766 27669 9818
rect 27693 9766 27723 9818
rect 27723 9766 27735 9818
rect 27735 9766 27749 9818
rect 27773 9766 27787 9818
rect 27787 9766 27799 9818
rect 27799 9766 27829 9818
rect 27853 9766 27863 9818
rect 27863 9766 27909 9818
rect 27613 9764 27669 9766
rect 27693 9764 27749 9766
rect 27773 9764 27829 9766
rect 27853 9764 27909 9766
rect 8178 9274 8234 9276
rect 8258 9274 8314 9276
rect 8338 9274 8394 9276
rect 8418 9274 8474 9276
rect 8178 9222 8224 9274
rect 8224 9222 8234 9274
rect 8258 9222 8288 9274
rect 8288 9222 8300 9274
rect 8300 9222 8314 9274
rect 8338 9222 8352 9274
rect 8352 9222 8364 9274
rect 8364 9222 8394 9274
rect 8418 9222 8428 9274
rect 8428 9222 8474 9274
rect 8178 9220 8234 9222
rect 8258 9220 8314 9222
rect 8338 9220 8394 9222
rect 8418 9220 8474 9222
rect 15952 9274 16008 9276
rect 16032 9274 16088 9276
rect 16112 9274 16168 9276
rect 16192 9274 16248 9276
rect 15952 9222 15998 9274
rect 15998 9222 16008 9274
rect 16032 9222 16062 9274
rect 16062 9222 16074 9274
rect 16074 9222 16088 9274
rect 16112 9222 16126 9274
rect 16126 9222 16138 9274
rect 16138 9222 16168 9274
rect 16192 9222 16202 9274
rect 16202 9222 16248 9274
rect 15952 9220 16008 9222
rect 16032 9220 16088 9222
rect 16112 9220 16168 9222
rect 16192 9220 16248 9222
rect 23726 9274 23782 9276
rect 23806 9274 23862 9276
rect 23886 9274 23942 9276
rect 23966 9274 24022 9276
rect 23726 9222 23772 9274
rect 23772 9222 23782 9274
rect 23806 9222 23836 9274
rect 23836 9222 23848 9274
rect 23848 9222 23862 9274
rect 23886 9222 23900 9274
rect 23900 9222 23912 9274
rect 23912 9222 23942 9274
rect 23966 9222 23976 9274
rect 23976 9222 24022 9274
rect 23726 9220 23782 9222
rect 23806 9220 23862 9222
rect 23886 9220 23942 9222
rect 23966 9220 24022 9222
rect 31500 9274 31556 9276
rect 31580 9274 31636 9276
rect 31660 9274 31716 9276
rect 31740 9274 31796 9276
rect 31500 9222 31546 9274
rect 31546 9222 31556 9274
rect 31580 9222 31610 9274
rect 31610 9222 31622 9274
rect 31622 9222 31636 9274
rect 31660 9222 31674 9274
rect 31674 9222 31686 9274
rect 31686 9222 31716 9274
rect 31740 9222 31750 9274
rect 31750 9222 31796 9274
rect 31500 9220 31556 9222
rect 31580 9220 31636 9222
rect 31660 9220 31716 9222
rect 31740 9220 31796 9222
rect 4291 8730 4347 8732
rect 4371 8730 4427 8732
rect 4451 8730 4507 8732
rect 4531 8730 4587 8732
rect 4291 8678 4337 8730
rect 4337 8678 4347 8730
rect 4371 8678 4401 8730
rect 4401 8678 4413 8730
rect 4413 8678 4427 8730
rect 4451 8678 4465 8730
rect 4465 8678 4477 8730
rect 4477 8678 4507 8730
rect 4531 8678 4541 8730
rect 4541 8678 4587 8730
rect 4291 8676 4347 8678
rect 4371 8676 4427 8678
rect 4451 8676 4507 8678
rect 4531 8676 4587 8678
rect 12065 8730 12121 8732
rect 12145 8730 12201 8732
rect 12225 8730 12281 8732
rect 12305 8730 12361 8732
rect 12065 8678 12111 8730
rect 12111 8678 12121 8730
rect 12145 8678 12175 8730
rect 12175 8678 12187 8730
rect 12187 8678 12201 8730
rect 12225 8678 12239 8730
rect 12239 8678 12251 8730
rect 12251 8678 12281 8730
rect 12305 8678 12315 8730
rect 12315 8678 12361 8730
rect 12065 8676 12121 8678
rect 12145 8676 12201 8678
rect 12225 8676 12281 8678
rect 12305 8676 12361 8678
rect 19839 8730 19895 8732
rect 19919 8730 19975 8732
rect 19999 8730 20055 8732
rect 20079 8730 20135 8732
rect 19839 8678 19885 8730
rect 19885 8678 19895 8730
rect 19919 8678 19949 8730
rect 19949 8678 19961 8730
rect 19961 8678 19975 8730
rect 19999 8678 20013 8730
rect 20013 8678 20025 8730
rect 20025 8678 20055 8730
rect 20079 8678 20089 8730
rect 20089 8678 20135 8730
rect 19839 8676 19895 8678
rect 19919 8676 19975 8678
rect 19999 8676 20055 8678
rect 20079 8676 20135 8678
rect 27613 8730 27669 8732
rect 27693 8730 27749 8732
rect 27773 8730 27829 8732
rect 27853 8730 27909 8732
rect 27613 8678 27659 8730
rect 27659 8678 27669 8730
rect 27693 8678 27723 8730
rect 27723 8678 27735 8730
rect 27735 8678 27749 8730
rect 27773 8678 27787 8730
rect 27787 8678 27799 8730
rect 27799 8678 27829 8730
rect 27853 8678 27863 8730
rect 27863 8678 27909 8730
rect 27613 8676 27669 8678
rect 27693 8676 27749 8678
rect 27773 8676 27829 8678
rect 27853 8676 27909 8678
rect 8178 8186 8234 8188
rect 8258 8186 8314 8188
rect 8338 8186 8394 8188
rect 8418 8186 8474 8188
rect 8178 8134 8224 8186
rect 8224 8134 8234 8186
rect 8258 8134 8288 8186
rect 8288 8134 8300 8186
rect 8300 8134 8314 8186
rect 8338 8134 8352 8186
rect 8352 8134 8364 8186
rect 8364 8134 8394 8186
rect 8418 8134 8428 8186
rect 8428 8134 8474 8186
rect 8178 8132 8234 8134
rect 8258 8132 8314 8134
rect 8338 8132 8394 8134
rect 8418 8132 8474 8134
rect 15952 8186 16008 8188
rect 16032 8186 16088 8188
rect 16112 8186 16168 8188
rect 16192 8186 16248 8188
rect 15952 8134 15998 8186
rect 15998 8134 16008 8186
rect 16032 8134 16062 8186
rect 16062 8134 16074 8186
rect 16074 8134 16088 8186
rect 16112 8134 16126 8186
rect 16126 8134 16138 8186
rect 16138 8134 16168 8186
rect 16192 8134 16202 8186
rect 16202 8134 16248 8186
rect 15952 8132 16008 8134
rect 16032 8132 16088 8134
rect 16112 8132 16168 8134
rect 16192 8132 16248 8134
rect 23726 8186 23782 8188
rect 23806 8186 23862 8188
rect 23886 8186 23942 8188
rect 23966 8186 24022 8188
rect 23726 8134 23772 8186
rect 23772 8134 23782 8186
rect 23806 8134 23836 8186
rect 23836 8134 23848 8186
rect 23848 8134 23862 8186
rect 23886 8134 23900 8186
rect 23900 8134 23912 8186
rect 23912 8134 23942 8186
rect 23966 8134 23976 8186
rect 23976 8134 24022 8186
rect 23726 8132 23782 8134
rect 23806 8132 23862 8134
rect 23886 8132 23942 8134
rect 23966 8132 24022 8134
rect 31500 8186 31556 8188
rect 31580 8186 31636 8188
rect 31660 8186 31716 8188
rect 31740 8186 31796 8188
rect 31500 8134 31546 8186
rect 31546 8134 31556 8186
rect 31580 8134 31610 8186
rect 31610 8134 31622 8186
rect 31622 8134 31636 8186
rect 31660 8134 31674 8186
rect 31674 8134 31686 8186
rect 31686 8134 31716 8186
rect 31740 8134 31750 8186
rect 31750 8134 31796 8186
rect 31500 8132 31556 8134
rect 31580 8132 31636 8134
rect 31660 8132 31716 8134
rect 31740 8132 31796 8134
rect 4291 7642 4347 7644
rect 4371 7642 4427 7644
rect 4451 7642 4507 7644
rect 4531 7642 4587 7644
rect 4291 7590 4337 7642
rect 4337 7590 4347 7642
rect 4371 7590 4401 7642
rect 4401 7590 4413 7642
rect 4413 7590 4427 7642
rect 4451 7590 4465 7642
rect 4465 7590 4477 7642
rect 4477 7590 4507 7642
rect 4531 7590 4541 7642
rect 4541 7590 4587 7642
rect 4291 7588 4347 7590
rect 4371 7588 4427 7590
rect 4451 7588 4507 7590
rect 4531 7588 4587 7590
rect 12065 7642 12121 7644
rect 12145 7642 12201 7644
rect 12225 7642 12281 7644
rect 12305 7642 12361 7644
rect 12065 7590 12111 7642
rect 12111 7590 12121 7642
rect 12145 7590 12175 7642
rect 12175 7590 12187 7642
rect 12187 7590 12201 7642
rect 12225 7590 12239 7642
rect 12239 7590 12251 7642
rect 12251 7590 12281 7642
rect 12305 7590 12315 7642
rect 12315 7590 12361 7642
rect 12065 7588 12121 7590
rect 12145 7588 12201 7590
rect 12225 7588 12281 7590
rect 12305 7588 12361 7590
rect 19839 7642 19895 7644
rect 19919 7642 19975 7644
rect 19999 7642 20055 7644
rect 20079 7642 20135 7644
rect 19839 7590 19885 7642
rect 19885 7590 19895 7642
rect 19919 7590 19949 7642
rect 19949 7590 19961 7642
rect 19961 7590 19975 7642
rect 19999 7590 20013 7642
rect 20013 7590 20025 7642
rect 20025 7590 20055 7642
rect 20079 7590 20089 7642
rect 20089 7590 20135 7642
rect 19839 7588 19895 7590
rect 19919 7588 19975 7590
rect 19999 7588 20055 7590
rect 20079 7588 20135 7590
rect 27613 7642 27669 7644
rect 27693 7642 27749 7644
rect 27773 7642 27829 7644
rect 27853 7642 27909 7644
rect 27613 7590 27659 7642
rect 27659 7590 27669 7642
rect 27693 7590 27723 7642
rect 27723 7590 27735 7642
rect 27735 7590 27749 7642
rect 27773 7590 27787 7642
rect 27787 7590 27799 7642
rect 27799 7590 27829 7642
rect 27853 7590 27863 7642
rect 27863 7590 27909 7642
rect 27613 7588 27669 7590
rect 27693 7588 27749 7590
rect 27773 7588 27829 7590
rect 27853 7588 27909 7590
rect 8178 7098 8234 7100
rect 8258 7098 8314 7100
rect 8338 7098 8394 7100
rect 8418 7098 8474 7100
rect 8178 7046 8224 7098
rect 8224 7046 8234 7098
rect 8258 7046 8288 7098
rect 8288 7046 8300 7098
rect 8300 7046 8314 7098
rect 8338 7046 8352 7098
rect 8352 7046 8364 7098
rect 8364 7046 8394 7098
rect 8418 7046 8428 7098
rect 8428 7046 8474 7098
rect 8178 7044 8234 7046
rect 8258 7044 8314 7046
rect 8338 7044 8394 7046
rect 8418 7044 8474 7046
rect 15952 7098 16008 7100
rect 16032 7098 16088 7100
rect 16112 7098 16168 7100
rect 16192 7098 16248 7100
rect 15952 7046 15998 7098
rect 15998 7046 16008 7098
rect 16032 7046 16062 7098
rect 16062 7046 16074 7098
rect 16074 7046 16088 7098
rect 16112 7046 16126 7098
rect 16126 7046 16138 7098
rect 16138 7046 16168 7098
rect 16192 7046 16202 7098
rect 16202 7046 16248 7098
rect 15952 7044 16008 7046
rect 16032 7044 16088 7046
rect 16112 7044 16168 7046
rect 16192 7044 16248 7046
rect 23726 7098 23782 7100
rect 23806 7098 23862 7100
rect 23886 7098 23942 7100
rect 23966 7098 24022 7100
rect 23726 7046 23772 7098
rect 23772 7046 23782 7098
rect 23806 7046 23836 7098
rect 23836 7046 23848 7098
rect 23848 7046 23862 7098
rect 23886 7046 23900 7098
rect 23900 7046 23912 7098
rect 23912 7046 23942 7098
rect 23966 7046 23976 7098
rect 23976 7046 24022 7098
rect 23726 7044 23782 7046
rect 23806 7044 23862 7046
rect 23886 7044 23942 7046
rect 23966 7044 24022 7046
rect 31500 7098 31556 7100
rect 31580 7098 31636 7100
rect 31660 7098 31716 7100
rect 31740 7098 31796 7100
rect 31500 7046 31546 7098
rect 31546 7046 31556 7098
rect 31580 7046 31610 7098
rect 31610 7046 31622 7098
rect 31622 7046 31636 7098
rect 31660 7046 31674 7098
rect 31674 7046 31686 7098
rect 31686 7046 31716 7098
rect 31740 7046 31750 7098
rect 31750 7046 31796 7098
rect 31500 7044 31556 7046
rect 31580 7044 31636 7046
rect 31660 7044 31716 7046
rect 31740 7044 31796 7046
rect 4291 6554 4347 6556
rect 4371 6554 4427 6556
rect 4451 6554 4507 6556
rect 4531 6554 4587 6556
rect 4291 6502 4337 6554
rect 4337 6502 4347 6554
rect 4371 6502 4401 6554
rect 4401 6502 4413 6554
rect 4413 6502 4427 6554
rect 4451 6502 4465 6554
rect 4465 6502 4477 6554
rect 4477 6502 4507 6554
rect 4531 6502 4541 6554
rect 4541 6502 4587 6554
rect 4291 6500 4347 6502
rect 4371 6500 4427 6502
rect 4451 6500 4507 6502
rect 4531 6500 4587 6502
rect 12065 6554 12121 6556
rect 12145 6554 12201 6556
rect 12225 6554 12281 6556
rect 12305 6554 12361 6556
rect 12065 6502 12111 6554
rect 12111 6502 12121 6554
rect 12145 6502 12175 6554
rect 12175 6502 12187 6554
rect 12187 6502 12201 6554
rect 12225 6502 12239 6554
rect 12239 6502 12251 6554
rect 12251 6502 12281 6554
rect 12305 6502 12315 6554
rect 12315 6502 12361 6554
rect 12065 6500 12121 6502
rect 12145 6500 12201 6502
rect 12225 6500 12281 6502
rect 12305 6500 12361 6502
rect 19839 6554 19895 6556
rect 19919 6554 19975 6556
rect 19999 6554 20055 6556
rect 20079 6554 20135 6556
rect 19839 6502 19885 6554
rect 19885 6502 19895 6554
rect 19919 6502 19949 6554
rect 19949 6502 19961 6554
rect 19961 6502 19975 6554
rect 19999 6502 20013 6554
rect 20013 6502 20025 6554
rect 20025 6502 20055 6554
rect 20079 6502 20089 6554
rect 20089 6502 20135 6554
rect 19839 6500 19895 6502
rect 19919 6500 19975 6502
rect 19999 6500 20055 6502
rect 20079 6500 20135 6502
rect 27613 6554 27669 6556
rect 27693 6554 27749 6556
rect 27773 6554 27829 6556
rect 27853 6554 27909 6556
rect 27613 6502 27659 6554
rect 27659 6502 27669 6554
rect 27693 6502 27723 6554
rect 27723 6502 27735 6554
rect 27735 6502 27749 6554
rect 27773 6502 27787 6554
rect 27787 6502 27799 6554
rect 27799 6502 27829 6554
rect 27853 6502 27863 6554
rect 27863 6502 27909 6554
rect 27613 6500 27669 6502
rect 27693 6500 27749 6502
rect 27773 6500 27829 6502
rect 27853 6500 27909 6502
rect 8178 6010 8234 6012
rect 8258 6010 8314 6012
rect 8338 6010 8394 6012
rect 8418 6010 8474 6012
rect 8178 5958 8224 6010
rect 8224 5958 8234 6010
rect 8258 5958 8288 6010
rect 8288 5958 8300 6010
rect 8300 5958 8314 6010
rect 8338 5958 8352 6010
rect 8352 5958 8364 6010
rect 8364 5958 8394 6010
rect 8418 5958 8428 6010
rect 8428 5958 8474 6010
rect 8178 5956 8234 5958
rect 8258 5956 8314 5958
rect 8338 5956 8394 5958
rect 8418 5956 8474 5958
rect 15952 6010 16008 6012
rect 16032 6010 16088 6012
rect 16112 6010 16168 6012
rect 16192 6010 16248 6012
rect 15952 5958 15998 6010
rect 15998 5958 16008 6010
rect 16032 5958 16062 6010
rect 16062 5958 16074 6010
rect 16074 5958 16088 6010
rect 16112 5958 16126 6010
rect 16126 5958 16138 6010
rect 16138 5958 16168 6010
rect 16192 5958 16202 6010
rect 16202 5958 16248 6010
rect 15952 5956 16008 5958
rect 16032 5956 16088 5958
rect 16112 5956 16168 5958
rect 16192 5956 16248 5958
rect 23726 6010 23782 6012
rect 23806 6010 23862 6012
rect 23886 6010 23942 6012
rect 23966 6010 24022 6012
rect 23726 5958 23772 6010
rect 23772 5958 23782 6010
rect 23806 5958 23836 6010
rect 23836 5958 23848 6010
rect 23848 5958 23862 6010
rect 23886 5958 23900 6010
rect 23900 5958 23912 6010
rect 23912 5958 23942 6010
rect 23966 5958 23976 6010
rect 23976 5958 24022 6010
rect 23726 5956 23782 5958
rect 23806 5956 23862 5958
rect 23886 5956 23942 5958
rect 23966 5956 24022 5958
rect 31500 6010 31556 6012
rect 31580 6010 31636 6012
rect 31660 6010 31716 6012
rect 31740 6010 31796 6012
rect 31500 5958 31546 6010
rect 31546 5958 31556 6010
rect 31580 5958 31610 6010
rect 31610 5958 31622 6010
rect 31622 5958 31636 6010
rect 31660 5958 31674 6010
rect 31674 5958 31686 6010
rect 31686 5958 31716 6010
rect 31740 5958 31750 6010
rect 31750 5958 31796 6010
rect 31500 5956 31556 5958
rect 31580 5956 31636 5958
rect 31660 5956 31716 5958
rect 31740 5956 31796 5958
rect 4291 5466 4347 5468
rect 4371 5466 4427 5468
rect 4451 5466 4507 5468
rect 4531 5466 4587 5468
rect 4291 5414 4337 5466
rect 4337 5414 4347 5466
rect 4371 5414 4401 5466
rect 4401 5414 4413 5466
rect 4413 5414 4427 5466
rect 4451 5414 4465 5466
rect 4465 5414 4477 5466
rect 4477 5414 4507 5466
rect 4531 5414 4541 5466
rect 4541 5414 4587 5466
rect 4291 5412 4347 5414
rect 4371 5412 4427 5414
rect 4451 5412 4507 5414
rect 4531 5412 4587 5414
rect 12065 5466 12121 5468
rect 12145 5466 12201 5468
rect 12225 5466 12281 5468
rect 12305 5466 12361 5468
rect 12065 5414 12111 5466
rect 12111 5414 12121 5466
rect 12145 5414 12175 5466
rect 12175 5414 12187 5466
rect 12187 5414 12201 5466
rect 12225 5414 12239 5466
rect 12239 5414 12251 5466
rect 12251 5414 12281 5466
rect 12305 5414 12315 5466
rect 12315 5414 12361 5466
rect 12065 5412 12121 5414
rect 12145 5412 12201 5414
rect 12225 5412 12281 5414
rect 12305 5412 12361 5414
rect 19839 5466 19895 5468
rect 19919 5466 19975 5468
rect 19999 5466 20055 5468
rect 20079 5466 20135 5468
rect 19839 5414 19885 5466
rect 19885 5414 19895 5466
rect 19919 5414 19949 5466
rect 19949 5414 19961 5466
rect 19961 5414 19975 5466
rect 19999 5414 20013 5466
rect 20013 5414 20025 5466
rect 20025 5414 20055 5466
rect 20079 5414 20089 5466
rect 20089 5414 20135 5466
rect 19839 5412 19895 5414
rect 19919 5412 19975 5414
rect 19999 5412 20055 5414
rect 20079 5412 20135 5414
rect 27613 5466 27669 5468
rect 27693 5466 27749 5468
rect 27773 5466 27829 5468
rect 27853 5466 27909 5468
rect 27613 5414 27659 5466
rect 27659 5414 27669 5466
rect 27693 5414 27723 5466
rect 27723 5414 27735 5466
rect 27735 5414 27749 5466
rect 27773 5414 27787 5466
rect 27787 5414 27799 5466
rect 27799 5414 27829 5466
rect 27853 5414 27863 5466
rect 27863 5414 27909 5466
rect 27613 5412 27669 5414
rect 27693 5412 27749 5414
rect 27773 5412 27829 5414
rect 27853 5412 27909 5414
rect 8178 4922 8234 4924
rect 8258 4922 8314 4924
rect 8338 4922 8394 4924
rect 8418 4922 8474 4924
rect 8178 4870 8224 4922
rect 8224 4870 8234 4922
rect 8258 4870 8288 4922
rect 8288 4870 8300 4922
rect 8300 4870 8314 4922
rect 8338 4870 8352 4922
rect 8352 4870 8364 4922
rect 8364 4870 8394 4922
rect 8418 4870 8428 4922
rect 8428 4870 8474 4922
rect 8178 4868 8234 4870
rect 8258 4868 8314 4870
rect 8338 4868 8394 4870
rect 8418 4868 8474 4870
rect 15952 4922 16008 4924
rect 16032 4922 16088 4924
rect 16112 4922 16168 4924
rect 16192 4922 16248 4924
rect 15952 4870 15998 4922
rect 15998 4870 16008 4922
rect 16032 4870 16062 4922
rect 16062 4870 16074 4922
rect 16074 4870 16088 4922
rect 16112 4870 16126 4922
rect 16126 4870 16138 4922
rect 16138 4870 16168 4922
rect 16192 4870 16202 4922
rect 16202 4870 16248 4922
rect 15952 4868 16008 4870
rect 16032 4868 16088 4870
rect 16112 4868 16168 4870
rect 16192 4868 16248 4870
rect 23726 4922 23782 4924
rect 23806 4922 23862 4924
rect 23886 4922 23942 4924
rect 23966 4922 24022 4924
rect 23726 4870 23772 4922
rect 23772 4870 23782 4922
rect 23806 4870 23836 4922
rect 23836 4870 23848 4922
rect 23848 4870 23862 4922
rect 23886 4870 23900 4922
rect 23900 4870 23912 4922
rect 23912 4870 23942 4922
rect 23966 4870 23976 4922
rect 23976 4870 24022 4922
rect 23726 4868 23782 4870
rect 23806 4868 23862 4870
rect 23886 4868 23942 4870
rect 23966 4868 24022 4870
rect 31500 4922 31556 4924
rect 31580 4922 31636 4924
rect 31660 4922 31716 4924
rect 31740 4922 31796 4924
rect 31500 4870 31546 4922
rect 31546 4870 31556 4922
rect 31580 4870 31610 4922
rect 31610 4870 31622 4922
rect 31622 4870 31636 4922
rect 31660 4870 31674 4922
rect 31674 4870 31686 4922
rect 31686 4870 31716 4922
rect 31740 4870 31750 4922
rect 31750 4870 31796 4922
rect 31500 4868 31556 4870
rect 31580 4868 31636 4870
rect 31660 4868 31716 4870
rect 31740 4868 31796 4870
rect 4291 4378 4347 4380
rect 4371 4378 4427 4380
rect 4451 4378 4507 4380
rect 4531 4378 4587 4380
rect 4291 4326 4337 4378
rect 4337 4326 4347 4378
rect 4371 4326 4401 4378
rect 4401 4326 4413 4378
rect 4413 4326 4427 4378
rect 4451 4326 4465 4378
rect 4465 4326 4477 4378
rect 4477 4326 4507 4378
rect 4531 4326 4541 4378
rect 4541 4326 4587 4378
rect 4291 4324 4347 4326
rect 4371 4324 4427 4326
rect 4451 4324 4507 4326
rect 4531 4324 4587 4326
rect 12065 4378 12121 4380
rect 12145 4378 12201 4380
rect 12225 4378 12281 4380
rect 12305 4378 12361 4380
rect 12065 4326 12111 4378
rect 12111 4326 12121 4378
rect 12145 4326 12175 4378
rect 12175 4326 12187 4378
rect 12187 4326 12201 4378
rect 12225 4326 12239 4378
rect 12239 4326 12251 4378
rect 12251 4326 12281 4378
rect 12305 4326 12315 4378
rect 12315 4326 12361 4378
rect 12065 4324 12121 4326
rect 12145 4324 12201 4326
rect 12225 4324 12281 4326
rect 12305 4324 12361 4326
rect 19839 4378 19895 4380
rect 19919 4378 19975 4380
rect 19999 4378 20055 4380
rect 20079 4378 20135 4380
rect 19839 4326 19885 4378
rect 19885 4326 19895 4378
rect 19919 4326 19949 4378
rect 19949 4326 19961 4378
rect 19961 4326 19975 4378
rect 19999 4326 20013 4378
rect 20013 4326 20025 4378
rect 20025 4326 20055 4378
rect 20079 4326 20089 4378
rect 20089 4326 20135 4378
rect 19839 4324 19895 4326
rect 19919 4324 19975 4326
rect 19999 4324 20055 4326
rect 20079 4324 20135 4326
rect 27613 4378 27669 4380
rect 27693 4378 27749 4380
rect 27773 4378 27829 4380
rect 27853 4378 27909 4380
rect 27613 4326 27659 4378
rect 27659 4326 27669 4378
rect 27693 4326 27723 4378
rect 27723 4326 27735 4378
rect 27735 4326 27749 4378
rect 27773 4326 27787 4378
rect 27787 4326 27799 4378
rect 27799 4326 27829 4378
rect 27853 4326 27863 4378
rect 27863 4326 27909 4378
rect 27613 4324 27669 4326
rect 27693 4324 27749 4326
rect 27773 4324 27829 4326
rect 27853 4324 27909 4326
rect 8178 3834 8234 3836
rect 8258 3834 8314 3836
rect 8338 3834 8394 3836
rect 8418 3834 8474 3836
rect 8178 3782 8224 3834
rect 8224 3782 8234 3834
rect 8258 3782 8288 3834
rect 8288 3782 8300 3834
rect 8300 3782 8314 3834
rect 8338 3782 8352 3834
rect 8352 3782 8364 3834
rect 8364 3782 8394 3834
rect 8418 3782 8428 3834
rect 8428 3782 8474 3834
rect 8178 3780 8234 3782
rect 8258 3780 8314 3782
rect 8338 3780 8394 3782
rect 8418 3780 8474 3782
rect 15952 3834 16008 3836
rect 16032 3834 16088 3836
rect 16112 3834 16168 3836
rect 16192 3834 16248 3836
rect 15952 3782 15998 3834
rect 15998 3782 16008 3834
rect 16032 3782 16062 3834
rect 16062 3782 16074 3834
rect 16074 3782 16088 3834
rect 16112 3782 16126 3834
rect 16126 3782 16138 3834
rect 16138 3782 16168 3834
rect 16192 3782 16202 3834
rect 16202 3782 16248 3834
rect 15952 3780 16008 3782
rect 16032 3780 16088 3782
rect 16112 3780 16168 3782
rect 16192 3780 16248 3782
rect 23726 3834 23782 3836
rect 23806 3834 23862 3836
rect 23886 3834 23942 3836
rect 23966 3834 24022 3836
rect 23726 3782 23772 3834
rect 23772 3782 23782 3834
rect 23806 3782 23836 3834
rect 23836 3782 23848 3834
rect 23848 3782 23862 3834
rect 23886 3782 23900 3834
rect 23900 3782 23912 3834
rect 23912 3782 23942 3834
rect 23966 3782 23976 3834
rect 23976 3782 24022 3834
rect 23726 3780 23782 3782
rect 23806 3780 23862 3782
rect 23886 3780 23942 3782
rect 23966 3780 24022 3782
rect 31500 3834 31556 3836
rect 31580 3834 31636 3836
rect 31660 3834 31716 3836
rect 31740 3834 31796 3836
rect 31500 3782 31546 3834
rect 31546 3782 31556 3834
rect 31580 3782 31610 3834
rect 31610 3782 31622 3834
rect 31622 3782 31636 3834
rect 31660 3782 31674 3834
rect 31674 3782 31686 3834
rect 31686 3782 31716 3834
rect 31740 3782 31750 3834
rect 31750 3782 31796 3834
rect 31500 3780 31556 3782
rect 31580 3780 31636 3782
rect 31660 3780 31716 3782
rect 31740 3780 31796 3782
rect 4291 3290 4347 3292
rect 4371 3290 4427 3292
rect 4451 3290 4507 3292
rect 4531 3290 4587 3292
rect 4291 3238 4337 3290
rect 4337 3238 4347 3290
rect 4371 3238 4401 3290
rect 4401 3238 4413 3290
rect 4413 3238 4427 3290
rect 4451 3238 4465 3290
rect 4465 3238 4477 3290
rect 4477 3238 4507 3290
rect 4531 3238 4541 3290
rect 4541 3238 4587 3290
rect 4291 3236 4347 3238
rect 4371 3236 4427 3238
rect 4451 3236 4507 3238
rect 4531 3236 4587 3238
rect 12065 3290 12121 3292
rect 12145 3290 12201 3292
rect 12225 3290 12281 3292
rect 12305 3290 12361 3292
rect 12065 3238 12111 3290
rect 12111 3238 12121 3290
rect 12145 3238 12175 3290
rect 12175 3238 12187 3290
rect 12187 3238 12201 3290
rect 12225 3238 12239 3290
rect 12239 3238 12251 3290
rect 12251 3238 12281 3290
rect 12305 3238 12315 3290
rect 12315 3238 12361 3290
rect 12065 3236 12121 3238
rect 12145 3236 12201 3238
rect 12225 3236 12281 3238
rect 12305 3236 12361 3238
rect 19839 3290 19895 3292
rect 19919 3290 19975 3292
rect 19999 3290 20055 3292
rect 20079 3290 20135 3292
rect 19839 3238 19885 3290
rect 19885 3238 19895 3290
rect 19919 3238 19949 3290
rect 19949 3238 19961 3290
rect 19961 3238 19975 3290
rect 19999 3238 20013 3290
rect 20013 3238 20025 3290
rect 20025 3238 20055 3290
rect 20079 3238 20089 3290
rect 20089 3238 20135 3290
rect 19839 3236 19895 3238
rect 19919 3236 19975 3238
rect 19999 3236 20055 3238
rect 20079 3236 20135 3238
rect 27613 3290 27669 3292
rect 27693 3290 27749 3292
rect 27773 3290 27829 3292
rect 27853 3290 27909 3292
rect 27613 3238 27659 3290
rect 27659 3238 27669 3290
rect 27693 3238 27723 3290
rect 27723 3238 27735 3290
rect 27735 3238 27749 3290
rect 27773 3238 27787 3290
rect 27787 3238 27799 3290
rect 27799 3238 27829 3290
rect 27853 3238 27863 3290
rect 27863 3238 27909 3290
rect 27613 3236 27669 3238
rect 27693 3236 27749 3238
rect 27773 3236 27829 3238
rect 27853 3236 27909 3238
rect 8178 2746 8234 2748
rect 8258 2746 8314 2748
rect 8338 2746 8394 2748
rect 8418 2746 8474 2748
rect 8178 2694 8224 2746
rect 8224 2694 8234 2746
rect 8258 2694 8288 2746
rect 8288 2694 8300 2746
rect 8300 2694 8314 2746
rect 8338 2694 8352 2746
rect 8352 2694 8364 2746
rect 8364 2694 8394 2746
rect 8418 2694 8428 2746
rect 8428 2694 8474 2746
rect 8178 2692 8234 2694
rect 8258 2692 8314 2694
rect 8338 2692 8394 2694
rect 8418 2692 8474 2694
rect 15952 2746 16008 2748
rect 16032 2746 16088 2748
rect 16112 2746 16168 2748
rect 16192 2746 16248 2748
rect 15952 2694 15998 2746
rect 15998 2694 16008 2746
rect 16032 2694 16062 2746
rect 16062 2694 16074 2746
rect 16074 2694 16088 2746
rect 16112 2694 16126 2746
rect 16126 2694 16138 2746
rect 16138 2694 16168 2746
rect 16192 2694 16202 2746
rect 16202 2694 16248 2746
rect 15952 2692 16008 2694
rect 16032 2692 16088 2694
rect 16112 2692 16168 2694
rect 16192 2692 16248 2694
rect 23726 2746 23782 2748
rect 23806 2746 23862 2748
rect 23886 2746 23942 2748
rect 23966 2746 24022 2748
rect 23726 2694 23772 2746
rect 23772 2694 23782 2746
rect 23806 2694 23836 2746
rect 23836 2694 23848 2746
rect 23848 2694 23862 2746
rect 23886 2694 23900 2746
rect 23900 2694 23912 2746
rect 23912 2694 23942 2746
rect 23966 2694 23976 2746
rect 23976 2694 24022 2746
rect 23726 2692 23782 2694
rect 23806 2692 23862 2694
rect 23886 2692 23942 2694
rect 23966 2692 24022 2694
rect 31500 2746 31556 2748
rect 31580 2746 31636 2748
rect 31660 2746 31716 2748
rect 31740 2746 31796 2748
rect 31500 2694 31546 2746
rect 31546 2694 31556 2746
rect 31580 2694 31610 2746
rect 31610 2694 31622 2746
rect 31622 2694 31636 2746
rect 31660 2694 31674 2746
rect 31674 2694 31686 2746
rect 31686 2694 31716 2746
rect 31740 2694 31750 2746
rect 31750 2694 31796 2746
rect 31500 2692 31556 2694
rect 31580 2692 31636 2694
rect 31660 2692 31716 2694
rect 31740 2692 31796 2694
rect 4291 2202 4347 2204
rect 4371 2202 4427 2204
rect 4451 2202 4507 2204
rect 4531 2202 4587 2204
rect 4291 2150 4337 2202
rect 4337 2150 4347 2202
rect 4371 2150 4401 2202
rect 4401 2150 4413 2202
rect 4413 2150 4427 2202
rect 4451 2150 4465 2202
rect 4465 2150 4477 2202
rect 4477 2150 4507 2202
rect 4531 2150 4541 2202
rect 4541 2150 4587 2202
rect 4291 2148 4347 2150
rect 4371 2148 4427 2150
rect 4451 2148 4507 2150
rect 4531 2148 4587 2150
rect 12065 2202 12121 2204
rect 12145 2202 12201 2204
rect 12225 2202 12281 2204
rect 12305 2202 12361 2204
rect 12065 2150 12111 2202
rect 12111 2150 12121 2202
rect 12145 2150 12175 2202
rect 12175 2150 12187 2202
rect 12187 2150 12201 2202
rect 12225 2150 12239 2202
rect 12239 2150 12251 2202
rect 12251 2150 12281 2202
rect 12305 2150 12315 2202
rect 12315 2150 12361 2202
rect 12065 2148 12121 2150
rect 12145 2148 12201 2150
rect 12225 2148 12281 2150
rect 12305 2148 12361 2150
rect 19839 2202 19895 2204
rect 19919 2202 19975 2204
rect 19999 2202 20055 2204
rect 20079 2202 20135 2204
rect 19839 2150 19885 2202
rect 19885 2150 19895 2202
rect 19919 2150 19949 2202
rect 19949 2150 19961 2202
rect 19961 2150 19975 2202
rect 19999 2150 20013 2202
rect 20013 2150 20025 2202
rect 20025 2150 20055 2202
rect 20079 2150 20089 2202
rect 20089 2150 20135 2202
rect 19839 2148 19895 2150
rect 19919 2148 19975 2150
rect 19999 2148 20055 2150
rect 20079 2148 20135 2150
rect 27613 2202 27669 2204
rect 27693 2202 27749 2204
rect 27773 2202 27829 2204
rect 27853 2202 27909 2204
rect 27613 2150 27659 2202
rect 27659 2150 27669 2202
rect 27693 2150 27723 2202
rect 27723 2150 27735 2202
rect 27735 2150 27749 2202
rect 27773 2150 27787 2202
rect 27787 2150 27799 2202
rect 27799 2150 27829 2202
rect 27853 2150 27863 2202
rect 27863 2150 27909 2202
rect 27613 2148 27669 2150
rect 27693 2148 27749 2150
rect 27773 2148 27829 2150
rect 27853 2148 27909 2150
rect 8178 1658 8234 1660
rect 8258 1658 8314 1660
rect 8338 1658 8394 1660
rect 8418 1658 8474 1660
rect 8178 1606 8224 1658
rect 8224 1606 8234 1658
rect 8258 1606 8288 1658
rect 8288 1606 8300 1658
rect 8300 1606 8314 1658
rect 8338 1606 8352 1658
rect 8352 1606 8364 1658
rect 8364 1606 8394 1658
rect 8418 1606 8428 1658
rect 8428 1606 8474 1658
rect 8178 1604 8234 1606
rect 8258 1604 8314 1606
rect 8338 1604 8394 1606
rect 8418 1604 8474 1606
rect 15952 1658 16008 1660
rect 16032 1658 16088 1660
rect 16112 1658 16168 1660
rect 16192 1658 16248 1660
rect 15952 1606 15998 1658
rect 15998 1606 16008 1658
rect 16032 1606 16062 1658
rect 16062 1606 16074 1658
rect 16074 1606 16088 1658
rect 16112 1606 16126 1658
rect 16126 1606 16138 1658
rect 16138 1606 16168 1658
rect 16192 1606 16202 1658
rect 16202 1606 16248 1658
rect 15952 1604 16008 1606
rect 16032 1604 16088 1606
rect 16112 1604 16168 1606
rect 16192 1604 16248 1606
rect 23726 1658 23782 1660
rect 23806 1658 23862 1660
rect 23886 1658 23942 1660
rect 23966 1658 24022 1660
rect 23726 1606 23772 1658
rect 23772 1606 23782 1658
rect 23806 1606 23836 1658
rect 23836 1606 23848 1658
rect 23848 1606 23862 1658
rect 23886 1606 23900 1658
rect 23900 1606 23912 1658
rect 23912 1606 23942 1658
rect 23966 1606 23976 1658
rect 23976 1606 24022 1658
rect 23726 1604 23782 1606
rect 23806 1604 23862 1606
rect 23886 1604 23942 1606
rect 23966 1604 24022 1606
rect 31500 1658 31556 1660
rect 31580 1658 31636 1660
rect 31660 1658 31716 1660
rect 31740 1658 31796 1660
rect 31500 1606 31546 1658
rect 31546 1606 31556 1658
rect 31580 1606 31610 1658
rect 31610 1606 31622 1658
rect 31622 1606 31636 1658
rect 31660 1606 31674 1658
rect 31674 1606 31686 1658
rect 31686 1606 31716 1658
rect 31740 1606 31750 1658
rect 31750 1606 31796 1658
rect 31500 1604 31556 1606
rect 31580 1604 31636 1606
rect 31660 1604 31716 1606
rect 31740 1604 31796 1606
rect 4291 1114 4347 1116
rect 4371 1114 4427 1116
rect 4451 1114 4507 1116
rect 4531 1114 4587 1116
rect 4291 1062 4337 1114
rect 4337 1062 4347 1114
rect 4371 1062 4401 1114
rect 4401 1062 4413 1114
rect 4413 1062 4427 1114
rect 4451 1062 4465 1114
rect 4465 1062 4477 1114
rect 4477 1062 4507 1114
rect 4531 1062 4541 1114
rect 4541 1062 4587 1114
rect 4291 1060 4347 1062
rect 4371 1060 4427 1062
rect 4451 1060 4507 1062
rect 4531 1060 4587 1062
rect 12065 1114 12121 1116
rect 12145 1114 12201 1116
rect 12225 1114 12281 1116
rect 12305 1114 12361 1116
rect 12065 1062 12111 1114
rect 12111 1062 12121 1114
rect 12145 1062 12175 1114
rect 12175 1062 12187 1114
rect 12187 1062 12201 1114
rect 12225 1062 12239 1114
rect 12239 1062 12251 1114
rect 12251 1062 12281 1114
rect 12305 1062 12315 1114
rect 12315 1062 12361 1114
rect 12065 1060 12121 1062
rect 12145 1060 12201 1062
rect 12225 1060 12281 1062
rect 12305 1060 12361 1062
rect 19839 1114 19895 1116
rect 19919 1114 19975 1116
rect 19999 1114 20055 1116
rect 20079 1114 20135 1116
rect 19839 1062 19885 1114
rect 19885 1062 19895 1114
rect 19919 1062 19949 1114
rect 19949 1062 19961 1114
rect 19961 1062 19975 1114
rect 19999 1062 20013 1114
rect 20013 1062 20025 1114
rect 20025 1062 20055 1114
rect 20079 1062 20089 1114
rect 20089 1062 20135 1114
rect 19839 1060 19895 1062
rect 19919 1060 19975 1062
rect 19999 1060 20055 1062
rect 20079 1060 20135 1062
rect 27613 1114 27669 1116
rect 27693 1114 27749 1116
rect 27773 1114 27829 1116
rect 27853 1114 27909 1116
rect 27613 1062 27659 1114
rect 27659 1062 27669 1114
rect 27693 1062 27723 1114
rect 27723 1062 27735 1114
rect 27735 1062 27749 1114
rect 27773 1062 27787 1114
rect 27787 1062 27799 1114
rect 27799 1062 27829 1114
rect 27853 1062 27863 1114
rect 27863 1062 27909 1114
rect 27613 1060 27669 1062
rect 27693 1060 27749 1062
rect 27773 1060 27829 1062
rect 27853 1060 27909 1062
rect 8178 570 8234 572
rect 8258 570 8314 572
rect 8338 570 8394 572
rect 8418 570 8474 572
rect 8178 518 8224 570
rect 8224 518 8234 570
rect 8258 518 8288 570
rect 8288 518 8300 570
rect 8300 518 8314 570
rect 8338 518 8352 570
rect 8352 518 8364 570
rect 8364 518 8394 570
rect 8418 518 8428 570
rect 8428 518 8474 570
rect 8178 516 8234 518
rect 8258 516 8314 518
rect 8338 516 8394 518
rect 8418 516 8474 518
rect 15952 570 16008 572
rect 16032 570 16088 572
rect 16112 570 16168 572
rect 16192 570 16248 572
rect 15952 518 15998 570
rect 15998 518 16008 570
rect 16032 518 16062 570
rect 16062 518 16074 570
rect 16074 518 16088 570
rect 16112 518 16126 570
rect 16126 518 16138 570
rect 16138 518 16168 570
rect 16192 518 16202 570
rect 16202 518 16248 570
rect 15952 516 16008 518
rect 16032 516 16088 518
rect 16112 516 16168 518
rect 16192 516 16248 518
rect 23726 570 23782 572
rect 23806 570 23862 572
rect 23886 570 23942 572
rect 23966 570 24022 572
rect 23726 518 23772 570
rect 23772 518 23782 570
rect 23806 518 23836 570
rect 23836 518 23848 570
rect 23848 518 23862 570
rect 23886 518 23900 570
rect 23900 518 23912 570
rect 23912 518 23942 570
rect 23966 518 23976 570
rect 23976 518 24022 570
rect 23726 516 23782 518
rect 23806 516 23862 518
rect 23886 516 23942 518
rect 23966 516 24022 518
rect 31500 570 31556 572
rect 31580 570 31636 572
rect 31660 570 31716 572
rect 31740 570 31796 572
rect 31500 518 31546 570
rect 31546 518 31556 570
rect 31580 518 31610 570
rect 31610 518 31622 570
rect 31622 518 31636 570
rect 31660 518 31674 570
rect 31674 518 31686 570
rect 31686 518 31716 570
rect 31740 518 31750 570
rect 31750 518 31796 570
rect 31500 516 31556 518
rect 31580 516 31636 518
rect 31660 516 31716 518
rect 31740 516 31796 518
<< metal3 >>
rect 28942 22266 28948 22268
rect 28820 22206 28948 22266
rect 28942 22204 28948 22206
rect 29012 22266 29018 22268
rect 29177 22266 29243 22269
rect 29012 22264 29243 22266
rect 29012 22208 29182 22264
rect 29238 22208 29243 22264
rect 29012 22206 29243 22208
rect 29012 22204 29018 22206
rect 29177 22203 29243 22206
rect 4521 21996 4587 21997
rect 4470 21932 4476 21996
rect 4540 21994 4587 21996
rect 4540 21992 4632 21994
rect 4582 21936 4632 21992
rect 4540 21934 4632 21936
rect 4540 21932 4587 21934
rect 8150 21932 8156 21996
rect 8220 21994 8226 21996
rect 8385 21994 8451 21997
rect 16297 21996 16363 21997
rect 8220 21992 8451 21994
rect 8220 21936 8390 21992
rect 8446 21936 8451 21992
rect 8220 21934 8451 21936
rect 8220 21932 8226 21934
rect 4521 21931 4587 21932
rect 8385 21931 8451 21934
rect 16246 21932 16252 21996
rect 16316 21994 16363 21996
rect 16316 21992 16408 21994
rect 16358 21936 16408 21992
rect 16316 21934 16408 21936
rect 16316 21932 16363 21934
rect 16297 21931 16363 21932
rect 841 21860 907 21861
rect 1577 21860 1643 21861
rect 2313 21860 2379 21861
rect 790 21796 796 21860
rect 860 21858 907 21860
rect 860 21856 952 21858
rect 902 21800 952 21856
rect 860 21798 952 21800
rect 860 21796 907 21798
rect 1526 21796 1532 21860
rect 1596 21858 1643 21860
rect 1596 21856 1688 21858
rect 1638 21800 1688 21856
rect 1596 21798 1688 21800
rect 1596 21796 1643 21798
rect 2262 21796 2268 21860
rect 2332 21858 2379 21860
rect 2332 21856 2424 21858
rect 2374 21800 2424 21856
rect 2332 21798 2424 21800
rect 2332 21796 2379 21798
rect 2998 21796 3004 21860
rect 3068 21858 3074 21860
rect 3233 21858 3299 21861
rect 3785 21860 3851 21861
rect 5257 21860 5323 21861
rect 5993 21860 6059 21861
rect 6729 21860 6795 21861
rect 7465 21860 7531 21861
rect 8937 21860 9003 21861
rect 9673 21860 9739 21861
rect 10409 21860 10475 21861
rect 11145 21860 11211 21861
rect 11881 21860 11947 21861
rect 12617 21860 12683 21861
rect 3068 21856 3299 21858
rect 3068 21800 3238 21856
rect 3294 21800 3299 21856
rect 3068 21798 3299 21800
rect 3068 21796 3074 21798
rect 841 21795 907 21796
rect 1577 21795 1643 21796
rect 2313 21795 2379 21796
rect 3233 21795 3299 21798
rect 3734 21796 3740 21860
rect 3804 21858 3851 21860
rect 3804 21856 3896 21858
rect 3846 21800 3896 21856
rect 3804 21798 3896 21800
rect 3804 21796 3851 21798
rect 5206 21796 5212 21860
rect 5276 21858 5323 21860
rect 5276 21856 5368 21858
rect 5318 21800 5368 21856
rect 5276 21798 5368 21800
rect 5276 21796 5323 21798
rect 5942 21796 5948 21860
rect 6012 21858 6059 21860
rect 6012 21856 6104 21858
rect 6054 21800 6104 21856
rect 6012 21798 6104 21800
rect 6012 21796 6059 21798
rect 6678 21796 6684 21860
rect 6748 21858 6795 21860
rect 6748 21856 6840 21858
rect 6790 21800 6840 21856
rect 6748 21798 6840 21800
rect 6748 21796 6795 21798
rect 7414 21796 7420 21860
rect 7484 21858 7531 21860
rect 7484 21856 7576 21858
rect 7526 21800 7576 21856
rect 7484 21798 7576 21800
rect 7484 21796 7531 21798
rect 8886 21796 8892 21860
rect 8956 21858 9003 21860
rect 8956 21856 9048 21858
rect 8998 21800 9048 21856
rect 8956 21798 9048 21800
rect 8956 21796 9003 21798
rect 9622 21796 9628 21860
rect 9692 21858 9739 21860
rect 9692 21856 9784 21858
rect 9734 21800 9784 21856
rect 9692 21798 9784 21800
rect 9692 21796 9739 21798
rect 10358 21796 10364 21860
rect 10428 21858 10475 21860
rect 10428 21856 10520 21858
rect 10470 21800 10520 21856
rect 10428 21798 10520 21800
rect 10428 21796 10475 21798
rect 11094 21796 11100 21860
rect 11164 21858 11211 21860
rect 11164 21856 11256 21858
rect 11206 21800 11256 21856
rect 11164 21798 11256 21800
rect 11164 21796 11211 21798
rect 11830 21796 11836 21860
rect 11900 21858 11947 21860
rect 11900 21856 11992 21858
rect 11942 21800 11992 21856
rect 11900 21798 11992 21800
rect 11900 21796 11947 21798
rect 12566 21796 12572 21860
rect 12636 21858 12683 21860
rect 12636 21856 12728 21858
rect 12678 21800 12728 21856
rect 12636 21798 12728 21800
rect 12636 21796 12683 21798
rect 13302 21796 13308 21860
rect 13372 21858 13378 21860
rect 13537 21858 13603 21861
rect 14089 21860 14155 21861
rect 14825 21860 14891 21861
rect 15561 21860 15627 21861
rect 17033 21860 17099 21861
rect 13372 21856 13603 21858
rect 13372 21800 13542 21856
rect 13598 21800 13603 21856
rect 13372 21798 13603 21800
rect 13372 21796 13378 21798
rect 3785 21795 3851 21796
rect 5257 21795 5323 21796
rect 5993 21795 6059 21796
rect 6729 21795 6795 21796
rect 7465 21795 7531 21796
rect 8937 21795 9003 21796
rect 9673 21795 9739 21796
rect 10409 21795 10475 21796
rect 11145 21795 11211 21796
rect 11881 21795 11947 21796
rect 12617 21795 12683 21796
rect 13537 21795 13603 21798
rect 14038 21796 14044 21860
rect 14108 21858 14155 21860
rect 14108 21856 14200 21858
rect 14150 21800 14200 21856
rect 14108 21798 14200 21800
rect 14108 21796 14155 21798
rect 14774 21796 14780 21860
rect 14844 21858 14891 21860
rect 14844 21856 14936 21858
rect 14886 21800 14936 21856
rect 14844 21798 14936 21800
rect 14844 21796 14891 21798
rect 15510 21796 15516 21860
rect 15580 21858 15627 21860
rect 15580 21856 15672 21858
rect 15622 21800 15672 21856
rect 15580 21798 15672 21800
rect 15580 21796 15627 21798
rect 16982 21796 16988 21860
rect 17052 21858 17099 21860
rect 17052 21856 17144 21858
rect 17094 21800 17144 21856
rect 17052 21798 17144 21800
rect 17052 21796 17099 21798
rect 29494 21796 29500 21860
rect 29564 21858 29570 21860
rect 29729 21858 29795 21861
rect 29564 21856 29795 21858
rect 29564 21800 29734 21856
rect 29790 21800 29795 21856
rect 29564 21798 29795 21800
rect 29564 21796 29570 21798
rect 14089 21795 14155 21796
rect 14825 21795 14891 21796
rect 15561 21795 15627 21796
rect 17033 21795 17099 21796
rect 29729 21795 29795 21798
rect 4281 21792 4597 21793
rect 4281 21728 4287 21792
rect 4351 21728 4367 21792
rect 4431 21728 4447 21792
rect 4511 21728 4527 21792
rect 4591 21728 4597 21792
rect 4281 21727 4597 21728
rect 12055 21792 12371 21793
rect 12055 21728 12061 21792
rect 12125 21728 12141 21792
rect 12205 21728 12221 21792
rect 12285 21728 12301 21792
rect 12365 21728 12371 21792
rect 12055 21727 12371 21728
rect 19829 21792 20145 21793
rect 19829 21728 19835 21792
rect 19899 21728 19915 21792
rect 19979 21728 19995 21792
rect 20059 21728 20075 21792
rect 20139 21728 20145 21792
rect 19829 21727 20145 21728
rect 27603 21792 27919 21793
rect 27603 21728 27609 21792
rect 27673 21728 27689 21792
rect 27753 21728 27769 21792
rect 27833 21728 27849 21792
rect 27913 21728 27919 21792
rect 27603 21727 27919 21728
rect 8168 21248 8484 21249
rect 8168 21184 8174 21248
rect 8238 21184 8254 21248
rect 8318 21184 8334 21248
rect 8398 21184 8414 21248
rect 8478 21184 8484 21248
rect 8168 21183 8484 21184
rect 15942 21248 16258 21249
rect 15942 21184 15948 21248
rect 16012 21184 16028 21248
rect 16092 21184 16108 21248
rect 16172 21184 16188 21248
rect 16252 21184 16258 21248
rect 15942 21183 16258 21184
rect 23716 21248 24032 21249
rect 23716 21184 23722 21248
rect 23786 21184 23802 21248
rect 23866 21184 23882 21248
rect 23946 21184 23962 21248
rect 24026 21184 24032 21248
rect 23716 21183 24032 21184
rect 31490 21248 31806 21249
rect 31490 21184 31496 21248
rect 31560 21184 31576 21248
rect 31640 21184 31656 21248
rect 31720 21184 31736 21248
rect 31800 21184 31806 21248
rect 31490 21183 31806 21184
rect 4281 20704 4597 20705
rect 4281 20640 4287 20704
rect 4351 20640 4367 20704
rect 4431 20640 4447 20704
rect 4511 20640 4527 20704
rect 4591 20640 4597 20704
rect 4281 20639 4597 20640
rect 12055 20704 12371 20705
rect 12055 20640 12061 20704
rect 12125 20640 12141 20704
rect 12205 20640 12221 20704
rect 12285 20640 12301 20704
rect 12365 20640 12371 20704
rect 12055 20639 12371 20640
rect 19829 20704 20145 20705
rect 19829 20640 19835 20704
rect 19899 20640 19915 20704
rect 19979 20640 19995 20704
rect 20059 20640 20075 20704
rect 20139 20640 20145 20704
rect 19829 20639 20145 20640
rect 27603 20704 27919 20705
rect 27603 20640 27609 20704
rect 27673 20640 27689 20704
rect 27753 20640 27769 20704
rect 27833 20640 27849 20704
rect 27913 20640 27919 20704
rect 27603 20639 27919 20640
rect 8168 20160 8484 20161
rect 8168 20096 8174 20160
rect 8238 20096 8254 20160
rect 8318 20096 8334 20160
rect 8398 20096 8414 20160
rect 8478 20096 8484 20160
rect 8168 20095 8484 20096
rect 15942 20160 16258 20161
rect 15942 20096 15948 20160
rect 16012 20096 16028 20160
rect 16092 20096 16108 20160
rect 16172 20096 16188 20160
rect 16252 20096 16258 20160
rect 15942 20095 16258 20096
rect 23716 20160 24032 20161
rect 23716 20096 23722 20160
rect 23786 20096 23802 20160
rect 23866 20096 23882 20160
rect 23946 20096 23962 20160
rect 24026 20096 24032 20160
rect 23716 20095 24032 20096
rect 31490 20160 31806 20161
rect 31490 20096 31496 20160
rect 31560 20096 31576 20160
rect 31640 20096 31656 20160
rect 31720 20096 31736 20160
rect 31800 20096 31806 20160
rect 31490 20095 31806 20096
rect 4281 19616 4597 19617
rect 4281 19552 4287 19616
rect 4351 19552 4367 19616
rect 4431 19552 4447 19616
rect 4511 19552 4527 19616
rect 4591 19552 4597 19616
rect 4281 19551 4597 19552
rect 12055 19616 12371 19617
rect 12055 19552 12061 19616
rect 12125 19552 12141 19616
rect 12205 19552 12221 19616
rect 12285 19552 12301 19616
rect 12365 19552 12371 19616
rect 12055 19551 12371 19552
rect 19829 19616 20145 19617
rect 19829 19552 19835 19616
rect 19899 19552 19915 19616
rect 19979 19552 19995 19616
rect 20059 19552 20075 19616
rect 20139 19552 20145 19616
rect 19829 19551 20145 19552
rect 27603 19616 27919 19617
rect 27603 19552 27609 19616
rect 27673 19552 27689 19616
rect 27753 19552 27769 19616
rect 27833 19552 27849 19616
rect 27913 19552 27919 19616
rect 27603 19551 27919 19552
rect 17718 19212 17724 19276
rect 17788 19274 17794 19276
rect 25681 19274 25747 19277
rect 17788 19272 25747 19274
rect 17788 19216 25686 19272
rect 25742 19216 25747 19272
rect 17788 19214 25747 19216
rect 17788 19212 17794 19214
rect 25681 19211 25747 19214
rect 8168 19072 8484 19073
rect 8168 19008 8174 19072
rect 8238 19008 8254 19072
rect 8318 19008 8334 19072
rect 8398 19008 8414 19072
rect 8478 19008 8484 19072
rect 8168 19007 8484 19008
rect 15942 19072 16258 19073
rect 15942 19008 15948 19072
rect 16012 19008 16028 19072
rect 16092 19008 16108 19072
rect 16172 19008 16188 19072
rect 16252 19008 16258 19072
rect 15942 19007 16258 19008
rect 23716 19072 24032 19073
rect 23716 19008 23722 19072
rect 23786 19008 23802 19072
rect 23866 19008 23882 19072
rect 23946 19008 23962 19072
rect 24026 19008 24032 19072
rect 23716 19007 24032 19008
rect 31490 19072 31806 19073
rect 31490 19008 31496 19072
rect 31560 19008 31576 19072
rect 31640 19008 31656 19072
rect 31720 19008 31736 19072
rect 31800 19008 31806 19072
rect 31490 19007 31806 19008
rect 4281 18528 4597 18529
rect 4281 18464 4287 18528
rect 4351 18464 4367 18528
rect 4431 18464 4447 18528
rect 4511 18464 4527 18528
rect 4591 18464 4597 18528
rect 4281 18463 4597 18464
rect 12055 18528 12371 18529
rect 12055 18464 12061 18528
rect 12125 18464 12141 18528
rect 12205 18464 12221 18528
rect 12285 18464 12301 18528
rect 12365 18464 12371 18528
rect 12055 18463 12371 18464
rect 19829 18528 20145 18529
rect 19829 18464 19835 18528
rect 19899 18464 19915 18528
rect 19979 18464 19995 18528
rect 20059 18464 20075 18528
rect 20139 18464 20145 18528
rect 19829 18463 20145 18464
rect 27603 18528 27919 18529
rect 27603 18464 27609 18528
rect 27673 18464 27689 18528
rect 27753 18464 27769 18528
rect 27833 18464 27849 18528
rect 27913 18464 27919 18528
rect 27603 18463 27919 18464
rect 8168 17984 8484 17985
rect 8168 17920 8174 17984
rect 8238 17920 8254 17984
rect 8318 17920 8334 17984
rect 8398 17920 8414 17984
rect 8478 17920 8484 17984
rect 8168 17919 8484 17920
rect 15942 17984 16258 17985
rect 15942 17920 15948 17984
rect 16012 17920 16028 17984
rect 16092 17920 16108 17984
rect 16172 17920 16188 17984
rect 16252 17920 16258 17984
rect 15942 17919 16258 17920
rect 23716 17984 24032 17985
rect 23716 17920 23722 17984
rect 23786 17920 23802 17984
rect 23866 17920 23882 17984
rect 23946 17920 23962 17984
rect 24026 17920 24032 17984
rect 23716 17919 24032 17920
rect 31490 17984 31806 17985
rect 31490 17920 31496 17984
rect 31560 17920 31576 17984
rect 31640 17920 31656 17984
rect 31720 17920 31736 17984
rect 31800 17920 31806 17984
rect 31490 17919 31806 17920
rect 4281 17440 4597 17441
rect 4281 17376 4287 17440
rect 4351 17376 4367 17440
rect 4431 17376 4447 17440
rect 4511 17376 4527 17440
rect 4591 17376 4597 17440
rect 4281 17375 4597 17376
rect 12055 17440 12371 17441
rect 12055 17376 12061 17440
rect 12125 17376 12141 17440
rect 12205 17376 12221 17440
rect 12285 17376 12301 17440
rect 12365 17376 12371 17440
rect 12055 17375 12371 17376
rect 19829 17440 20145 17441
rect 19829 17376 19835 17440
rect 19899 17376 19915 17440
rect 19979 17376 19995 17440
rect 20059 17376 20075 17440
rect 20139 17376 20145 17440
rect 19829 17375 20145 17376
rect 27603 17440 27919 17441
rect 27603 17376 27609 17440
rect 27673 17376 27689 17440
rect 27753 17376 27769 17440
rect 27833 17376 27849 17440
rect 27913 17376 27919 17440
rect 27603 17375 27919 17376
rect 8168 16896 8484 16897
rect 8168 16832 8174 16896
rect 8238 16832 8254 16896
rect 8318 16832 8334 16896
rect 8398 16832 8414 16896
rect 8478 16832 8484 16896
rect 8168 16831 8484 16832
rect 15942 16896 16258 16897
rect 15942 16832 15948 16896
rect 16012 16832 16028 16896
rect 16092 16832 16108 16896
rect 16172 16832 16188 16896
rect 16252 16832 16258 16896
rect 15942 16831 16258 16832
rect 23716 16896 24032 16897
rect 23716 16832 23722 16896
rect 23786 16832 23802 16896
rect 23866 16832 23882 16896
rect 23946 16832 23962 16896
rect 24026 16832 24032 16896
rect 23716 16831 24032 16832
rect 31490 16896 31806 16897
rect 31490 16832 31496 16896
rect 31560 16832 31576 16896
rect 31640 16832 31656 16896
rect 31720 16832 31736 16896
rect 31800 16832 31806 16896
rect 31490 16831 31806 16832
rect 4281 16352 4597 16353
rect 4281 16288 4287 16352
rect 4351 16288 4367 16352
rect 4431 16288 4447 16352
rect 4511 16288 4527 16352
rect 4591 16288 4597 16352
rect 4281 16287 4597 16288
rect 12055 16352 12371 16353
rect 12055 16288 12061 16352
rect 12125 16288 12141 16352
rect 12205 16288 12221 16352
rect 12285 16288 12301 16352
rect 12365 16288 12371 16352
rect 12055 16287 12371 16288
rect 19829 16352 20145 16353
rect 19829 16288 19835 16352
rect 19899 16288 19915 16352
rect 19979 16288 19995 16352
rect 20059 16288 20075 16352
rect 20139 16288 20145 16352
rect 19829 16287 20145 16288
rect 27603 16352 27919 16353
rect 27603 16288 27609 16352
rect 27673 16288 27689 16352
rect 27753 16288 27769 16352
rect 27833 16288 27849 16352
rect 27913 16288 27919 16352
rect 27603 16287 27919 16288
rect 8168 15808 8484 15809
rect 8168 15744 8174 15808
rect 8238 15744 8254 15808
rect 8318 15744 8334 15808
rect 8398 15744 8414 15808
rect 8478 15744 8484 15808
rect 8168 15743 8484 15744
rect 15942 15808 16258 15809
rect 15942 15744 15948 15808
rect 16012 15744 16028 15808
rect 16092 15744 16108 15808
rect 16172 15744 16188 15808
rect 16252 15744 16258 15808
rect 15942 15743 16258 15744
rect 23716 15808 24032 15809
rect 23716 15744 23722 15808
rect 23786 15744 23802 15808
rect 23866 15744 23882 15808
rect 23946 15744 23962 15808
rect 24026 15744 24032 15808
rect 23716 15743 24032 15744
rect 31490 15808 31806 15809
rect 31490 15744 31496 15808
rect 31560 15744 31576 15808
rect 31640 15744 31656 15808
rect 31720 15744 31736 15808
rect 31800 15744 31806 15808
rect 31490 15743 31806 15744
rect 4281 15264 4597 15265
rect 4281 15200 4287 15264
rect 4351 15200 4367 15264
rect 4431 15200 4447 15264
rect 4511 15200 4527 15264
rect 4591 15200 4597 15264
rect 4281 15199 4597 15200
rect 12055 15264 12371 15265
rect 12055 15200 12061 15264
rect 12125 15200 12141 15264
rect 12205 15200 12221 15264
rect 12285 15200 12301 15264
rect 12365 15200 12371 15264
rect 12055 15199 12371 15200
rect 19829 15264 20145 15265
rect 19829 15200 19835 15264
rect 19899 15200 19915 15264
rect 19979 15200 19995 15264
rect 20059 15200 20075 15264
rect 20139 15200 20145 15264
rect 19829 15199 20145 15200
rect 27603 15264 27919 15265
rect 27603 15200 27609 15264
rect 27673 15200 27689 15264
rect 27753 15200 27769 15264
rect 27833 15200 27849 15264
rect 27913 15200 27919 15264
rect 27603 15199 27919 15200
rect 8168 14720 8484 14721
rect 8168 14656 8174 14720
rect 8238 14656 8254 14720
rect 8318 14656 8334 14720
rect 8398 14656 8414 14720
rect 8478 14656 8484 14720
rect 8168 14655 8484 14656
rect 15942 14720 16258 14721
rect 15942 14656 15948 14720
rect 16012 14656 16028 14720
rect 16092 14656 16108 14720
rect 16172 14656 16188 14720
rect 16252 14656 16258 14720
rect 15942 14655 16258 14656
rect 23716 14720 24032 14721
rect 23716 14656 23722 14720
rect 23786 14656 23802 14720
rect 23866 14656 23882 14720
rect 23946 14656 23962 14720
rect 24026 14656 24032 14720
rect 23716 14655 24032 14656
rect 31490 14720 31806 14721
rect 31490 14656 31496 14720
rect 31560 14656 31576 14720
rect 31640 14656 31656 14720
rect 31720 14656 31736 14720
rect 31800 14656 31806 14720
rect 31490 14655 31806 14656
rect 4281 14176 4597 14177
rect 4281 14112 4287 14176
rect 4351 14112 4367 14176
rect 4431 14112 4447 14176
rect 4511 14112 4527 14176
rect 4591 14112 4597 14176
rect 4281 14111 4597 14112
rect 12055 14176 12371 14177
rect 12055 14112 12061 14176
rect 12125 14112 12141 14176
rect 12205 14112 12221 14176
rect 12285 14112 12301 14176
rect 12365 14112 12371 14176
rect 12055 14111 12371 14112
rect 19829 14176 20145 14177
rect 19829 14112 19835 14176
rect 19899 14112 19915 14176
rect 19979 14112 19995 14176
rect 20059 14112 20075 14176
rect 20139 14112 20145 14176
rect 19829 14111 20145 14112
rect 27603 14176 27919 14177
rect 27603 14112 27609 14176
rect 27673 14112 27689 14176
rect 27753 14112 27769 14176
rect 27833 14112 27849 14176
rect 27913 14112 27919 14176
rect 27603 14111 27919 14112
rect 8168 13632 8484 13633
rect 8168 13568 8174 13632
rect 8238 13568 8254 13632
rect 8318 13568 8334 13632
rect 8398 13568 8414 13632
rect 8478 13568 8484 13632
rect 8168 13567 8484 13568
rect 15942 13632 16258 13633
rect 15942 13568 15948 13632
rect 16012 13568 16028 13632
rect 16092 13568 16108 13632
rect 16172 13568 16188 13632
rect 16252 13568 16258 13632
rect 15942 13567 16258 13568
rect 23716 13632 24032 13633
rect 23716 13568 23722 13632
rect 23786 13568 23802 13632
rect 23866 13568 23882 13632
rect 23946 13568 23962 13632
rect 24026 13568 24032 13632
rect 23716 13567 24032 13568
rect 31490 13632 31806 13633
rect 31490 13568 31496 13632
rect 31560 13568 31576 13632
rect 31640 13568 31656 13632
rect 31720 13568 31736 13632
rect 31800 13568 31806 13632
rect 31490 13567 31806 13568
rect 4281 13088 4597 13089
rect 4281 13024 4287 13088
rect 4351 13024 4367 13088
rect 4431 13024 4447 13088
rect 4511 13024 4527 13088
rect 4591 13024 4597 13088
rect 4281 13023 4597 13024
rect 12055 13088 12371 13089
rect 12055 13024 12061 13088
rect 12125 13024 12141 13088
rect 12205 13024 12221 13088
rect 12285 13024 12301 13088
rect 12365 13024 12371 13088
rect 12055 13023 12371 13024
rect 19829 13088 20145 13089
rect 19829 13024 19835 13088
rect 19899 13024 19915 13088
rect 19979 13024 19995 13088
rect 20059 13024 20075 13088
rect 20139 13024 20145 13088
rect 19829 13023 20145 13024
rect 27603 13088 27919 13089
rect 27603 13024 27609 13088
rect 27673 13024 27689 13088
rect 27753 13024 27769 13088
rect 27833 13024 27849 13088
rect 27913 13024 27919 13088
rect 27603 13023 27919 13024
rect 8168 12544 8484 12545
rect 8168 12480 8174 12544
rect 8238 12480 8254 12544
rect 8318 12480 8334 12544
rect 8398 12480 8414 12544
rect 8478 12480 8484 12544
rect 8168 12479 8484 12480
rect 15942 12544 16258 12545
rect 15942 12480 15948 12544
rect 16012 12480 16028 12544
rect 16092 12480 16108 12544
rect 16172 12480 16188 12544
rect 16252 12480 16258 12544
rect 15942 12479 16258 12480
rect 23716 12544 24032 12545
rect 23716 12480 23722 12544
rect 23786 12480 23802 12544
rect 23866 12480 23882 12544
rect 23946 12480 23962 12544
rect 24026 12480 24032 12544
rect 23716 12479 24032 12480
rect 31490 12544 31806 12545
rect 31490 12480 31496 12544
rect 31560 12480 31576 12544
rect 31640 12480 31656 12544
rect 31720 12480 31736 12544
rect 31800 12480 31806 12544
rect 31490 12479 31806 12480
rect 4281 12000 4597 12001
rect 4281 11936 4287 12000
rect 4351 11936 4367 12000
rect 4431 11936 4447 12000
rect 4511 11936 4527 12000
rect 4591 11936 4597 12000
rect 4281 11935 4597 11936
rect 12055 12000 12371 12001
rect 12055 11936 12061 12000
rect 12125 11936 12141 12000
rect 12205 11936 12221 12000
rect 12285 11936 12301 12000
rect 12365 11936 12371 12000
rect 12055 11935 12371 11936
rect 19829 12000 20145 12001
rect 19829 11936 19835 12000
rect 19899 11936 19915 12000
rect 19979 11936 19995 12000
rect 20059 11936 20075 12000
rect 20139 11936 20145 12000
rect 19829 11935 20145 11936
rect 27603 12000 27919 12001
rect 27603 11936 27609 12000
rect 27673 11936 27689 12000
rect 27753 11936 27769 12000
rect 27833 11936 27849 12000
rect 27913 11936 27919 12000
rect 27603 11935 27919 11936
rect 8168 11456 8484 11457
rect 8168 11392 8174 11456
rect 8238 11392 8254 11456
rect 8318 11392 8334 11456
rect 8398 11392 8414 11456
rect 8478 11392 8484 11456
rect 8168 11391 8484 11392
rect 15942 11456 16258 11457
rect 15942 11392 15948 11456
rect 16012 11392 16028 11456
rect 16092 11392 16108 11456
rect 16172 11392 16188 11456
rect 16252 11392 16258 11456
rect 15942 11391 16258 11392
rect 23716 11456 24032 11457
rect 23716 11392 23722 11456
rect 23786 11392 23802 11456
rect 23866 11392 23882 11456
rect 23946 11392 23962 11456
rect 24026 11392 24032 11456
rect 23716 11391 24032 11392
rect 31490 11456 31806 11457
rect 31490 11392 31496 11456
rect 31560 11392 31576 11456
rect 31640 11392 31656 11456
rect 31720 11392 31736 11456
rect 31800 11392 31806 11456
rect 31490 11391 31806 11392
rect 4281 10912 4597 10913
rect 4281 10848 4287 10912
rect 4351 10848 4367 10912
rect 4431 10848 4447 10912
rect 4511 10848 4527 10912
rect 4591 10848 4597 10912
rect 4281 10847 4597 10848
rect 12055 10912 12371 10913
rect 12055 10848 12061 10912
rect 12125 10848 12141 10912
rect 12205 10848 12221 10912
rect 12285 10848 12301 10912
rect 12365 10848 12371 10912
rect 12055 10847 12371 10848
rect 19829 10912 20145 10913
rect 19829 10848 19835 10912
rect 19899 10848 19915 10912
rect 19979 10848 19995 10912
rect 20059 10848 20075 10912
rect 20139 10848 20145 10912
rect 19829 10847 20145 10848
rect 27603 10912 27919 10913
rect 27603 10848 27609 10912
rect 27673 10848 27689 10912
rect 27753 10848 27769 10912
rect 27833 10848 27849 10912
rect 27913 10848 27919 10912
rect 27603 10847 27919 10848
rect 8168 10368 8484 10369
rect 8168 10304 8174 10368
rect 8238 10304 8254 10368
rect 8318 10304 8334 10368
rect 8398 10304 8414 10368
rect 8478 10304 8484 10368
rect 8168 10303 8484 10304
rect 15942 10368 16258 10369
rect 15942 10304 15948 10368
rect 16012 10304 16028 10368
rect 16092 10304 16108 10368
rect 16172 10304 16188 10368
rect 16252 10304 16258 10368
rect 15942 10303 16258 10304
rect 23716 10368 24032 10369
rect 23716 10304 23722 10368
rect 23786 10304 23802 10368
rect 23866 10304 23882 10368
rect 23946 10304 23962 10368
rect 24026 10304 24032 10368
rect 23716 10303 24032 10304
rect 31490 10368 31806 10369
rect 31490 10304 31496 10368
rect 31560 10304 31576 10368
rect 31640 10304 31656 10368
rect 31720 10304 31736 10368
rect 31800 10304 31806 10368
rect 31490 10303 31806 10304
rect 4281 9824 4597 9825
rect 4281 9760 4287 9824
rect 4351 9760 4367 9824
rect 4431 9760 4447 9824
rect 4511 9760 4527 9824
rect 4591 9760 4597 9824
rect 4281 9759 4597 9760
rect 12055 9824 12371 9825
rect 12055 9760 12061 9824
rect 12125 9760 12141 9824
rect 12205 9760 12221 9824
rect 12285 9760 12301 9824
rect 12365 9760 12371 9824
rect 12055 9759 12371 9760
rect 19829 9824 20145 9825
rect 19829 9760 19835 9824
rect 19899 9760 19915 9824
rect 19979 9760 19995 9824
rect 20059 9760 20075 9824
rect 20139 9760 20145 9824
rect 19829 9759 20145 9760
rect 27603 9824 27919 9825
rect 27603 9760 27609 9824
rect 27673 9760 27689 9824
rect 27753 9760 27769 9824
rect 27833 9760 27849 9824
rect 27913 9760 27919 9824
rect 27603 9759 27919 9760
rect 8168 9280 8484 9281
rect 8168 9216 8174 9280
rect 8238 9216 8254 9280
rect 8318 9216 8334 9280
rect 8398 9216 8414 9280
rect 8478 9216 8484 9280
rect 8168 9215 8484 9216
rect 15942 9280 16258 9281
rect 15942 9216 15948 9280
rect 16012 9216 16028 9280
rect 16092 9216 16108 9280
rect 16172 9216 16188 9280
rect 16252 9216 16258 9280
rect 15942 9215 16258 9216
rect 23716 9280 24032 9281
rect 23716 9216 23722 9280
rect 23786 9216 23802 9280
rect 23866 9216 23882 9280
rect 23946 9216 23962 9280
rect 24026 9216 24032 9280
rect 23716 9215 24032 9216
rect 31490 9280 31806 9281
rect 31490 9216 31496 9280
rect 31560 9216 31576 9280
rect 31640 9216 31656 9280
rect 31720 9216 31736 9280
rect 31800 9216 31806 9280
rect 31490 9215 31806 9216
rect 4281 8736 4597 8737
rect 4281 8672 4287 8736
rect 4351 8672 4367 8736
rect 4431 8672 4447 8736
rect 4511 8672 4527 8736
rect 4591 8672 4597 8736
rect 4281 8671 4597 8672
rect 12055 8736 12371 8737
rect 12055 8672 12061 8736
rect 12125 8672 12141 8736
rect 12205 8672 12221 8736
rect 12285 8672 12301 8736
rect 12365 8672 12371 8736
rect 12055 8671 12371 8672
rect 19829 8736 20145 8737
rect 19829 8672 19835 8736
rect 19899 8672 19915 8736
rect 19979 8672 19995 8736
rect 20059 8672 20075 8736
rect 20139 8672 20145 8736
rect 19829 8671 20145 8672
rect 27603 8736 27919 8737
rect 27603 8672 27609 8736
rect 27673 8672 27689 8736
rect 27753 8672 27769 8736
rect 27833 8672 27849 8736
rect 27913 8672 27919 8736
rect 27603 8671 27919 8672
rect 8168 8192 8484 8193
rect 8168 8128 8174 8192
rect 8238 8128 8254 8192
rect 8318 8128 8334 8192
rect 8398 8128 8414 8192
rect 8478 8128 8484 8192
rect 8168 8127 8484 8128
rect 15942 8192 16258 8193
rect 15942 8128 15948 8192
rect 16012 8128 16028 8192
rect 16092 8128 16108 8192
rect 16172 8128 16188 8192
rect 16252 8128 16258 8192
rect 15942 8127 16258 8128
rect 23716 8192 24032 8193
rect 23716 8128 23722 8192
rect 23786 8128 23802 8192
rect 23866 8128 23882 8192
rect 23946 8128 23962 8192
rect 24026 8128 24032 8192
rect 23716 8127 24032 8128
rect 31490 8192 31806 8193
rect 31490 8128 31496 8192
rect 31560 8128 31576 8192
rect 31640 8128 31656 8192
rect 31720 8128 31736 8192
rect 31800 8128 31806 8192
rect 31490 8127 31806 8128
rect 4281 7648 4597 7649
rect 4281 7584 4287 7648
rect 4351 7584 4367 7648
rect 4431 7584 4447 7648
rect 4511 7584 4527 7648
rect 4591 7584 4597 7648
rect 4281 7583 4597 7584
rect 12055 7648 12371 7649
rect 12055 7584 12061 7648
rect 12125 7584 12141 7648
rect 12205 7584 12221 7648
rect 12285 7584 12301 7648
rect 12365 7584 12371 7648
rect 12055 7583 12371 7584
rect 19829 7648 20145 7649
rect 19829 7584 19835 7648
rect 19899 7584 19915 7648
rect 19979 7584 19995 7648
rect 20059 7584 20075 7648
rect 20139 7584 20145 7648
rect 19829 7583 20145 7584
rect 27603 7648 27919 7649
rect 27603 7584 27609 7648
rect 27673 7584 27689 7648
rect 27753 7584 27769 7648
rect 27833 7584 27849 7648
rect 27913 7584 27919 7648
rect 27603 7583 27919 7584
rect 8168 7104 8484 7105
rect 8168 7040 8174 7104
rect 8238 7040 8254 7104
rect 8318 7040 8334 7104
rect 8398 7040 8414 7104
rect 8478 7040 8484 7104
rect 8168 7039 8484 7040
rect 15942 7104 16258 7105
rect 15942 7040 15948 7104
rect 16012 7040 16028 7104
rect 16092 7040 16108 7104
rect 16172 7040 16188 7104
rect 16252 7040 16258 7104
rect 15942 7039 16258 7040
rect 23716 7104 24032 7105
rect 23716 7040 23722 7104
rect 23786 7040 23802 7104
rect 23866 7040 23882 7104
rect 23946 7040 23962 7104
rect 24026 7040 24032 7104
rect 23716 7039 24032 7040
rect 31490 7104 31806 7105
rect 31490 7040 31496 7104
rect 31560 7040 31576 7104
rect 31640 7040 31656 7104
rect 31720 7040 31736 7104
rect 31800 7040 31806 7104
rect 31490 7039 31806 7040
rect 4281 6560 4597 6561
rect 4281 6496 4287 6560
rect 4351 6496 4367 6560
rect 4431 6496 4447 6560
rect 4511 6496 4527 6560
rect 4591 6496 4597 6560
rect 4281 6495 4597 6496
rect 12055 6560 12371 6561
rect 12055 6496 12061 6560
rect 12125 6496 12141 6560
rect 12205 6496 12221 6560
rect 12285 6496 12301 6560
rect 12365 6496 12371 6560
rect 12055 6495 12371 6496
rect 19829 6560 20145 6561
rect 19829 6496 19835 6560
rect 19899 6496 19915 6560
rect 19979 6496 19995 6560
rect 20059 6496 20075 6560
rect 20139 6496 20145 6560
rect 19829 6495 20145 6496
rect 27603 6560 27919 6561
rect 27603 6496 27609 6560
rect 27673 6496 27689 6560
rect 27753 6496 27769 6560
rect 27833 6496 27849 6560
rect 27913 6496 27919 6560
rect 27603 6495 27919 6496
rect 8168 6016 8484 6017
rect 8168 5952 8174 6016
rect 8238 5952 8254 6016
rect 8318 5952 8334 6016
rect 8398 5952 8414 6016
rect 8478 5952 8484 6016
rect 8168 5951 8484 5952
rect 15942 6016 16258 6017
rect 15942 5952 15948 6016
rect 16012 5952 16028 6016
rect 16092 5952 16108 6016
rect 16172 5952 16188 6016
rect 16252 5952 16258 6016
rect 15942 5951 16258 5952
rect 23716 6016 24032 6017
rect 23716 5952 23722 6016
rect 23786 5952 23802 6016
rect 23866 5952 23882 6016
rect 23946 5952 23962 6016
rect 24026 5952 24032 6016
rect 23716 5951 24032 5952
rect 31490 6016 31806 6017
rect 31490 5952 31496 6016
rect 31560 5952 31576 6016
rect 31640 5952 31656 6016
rect 31720 5952 31736 6016
rect 31800 5952 31806 6016
rect 31490 5951 31806 5952
rect 4281 5472 4597 5473
rect 4281 5408 4287 5472
rect 4351 5408 4367 5472
rect 4431 5408 4447 5472
rect 4511 5408 4527 5472
rect 4591 5408 4597 5472
rect 4281 5407 4597 5408
rect 12055 5472 12371 5473
rect 12055 5408 12061 5472
rect 12125 5408 12141 5472
rect 12205 5408 12221 5472
rect 12285 5408 12301 5472
rect 12365 5408 12371 5472
rect 12055 5407 12371 5408
rect 19829 5472 20145 5473
rect 19829 5408 19835 5472
rect 19899 5408 19915 5472
rect 19979 5408 19995 5472
rect 20059 5408 20075 5472
rect 20139 5408 20145 5472
rect 19829 5407 20145 5408
rect 27603 5472 27919 5473
rect 27603 5408 27609 5472
rect 27673 5408 27689 5472
rect 27753 5408 27769 5472
rect 27833 5408 27849 5472
rect 27913 5408 27919 5472
rect 27603 5407 27919 5408
rect 8168 4928 8484 4929
rect 8168 4864 8174 4928
rect 8238 4864 8254 4928
rect 8318 4864 8334 4928
rect 8398 4864 8414 4928
rect 8478 4864 8484 4928
rect 8168 4863 8484 4864
rect 15942 4928 16258 4929
rect 15942 4864 15948 4928
rect 16012 4864 16028 4928
rect 16092 4864 16108 4928
rect 16172 4864 16188 4928
rect 16252 4864 16258 4928
rect 15942 4863 16258 4864
rect 23716 4928 24032 4929
rect 23716 4864 23722 4928
rect 23786 4864 23802 4928
rect 23866 4864 23882 4928
rect 23946 4864 23962 4928
rect 24026 4864 24032 4928
rect 23716 4863 24032 4864
rect 31490 4928 31806 4929
rect 31490 4864 31496 4928
rect 31560 4864 31576 4928
rect 31640 4864 31656 4928
rect 31720 4864 31736 4928
rect 31800 4864 31806 4928
rect 31490 4863 31806 4864
rect 4281 4384 4597 4385
rect 4281 4320 4287 4384
rect 4351 4320 4367 4384
rect 4431 4320 4447 4384
rect 4511 4320 4527 4384
rect 4591 4320 4597 4384
rect 4281 4319 4597 4320
rect 12055 4384 12371 4385
rect 12055 4320 12061 4384
rect 12125 4320 12141 4384
rect 12205 4320 12221 4384
rect 12285 4320 12301 4384
rect 12365 4320 12371 4384
rect 12055 4319 12371 4320
rect 19829 4384 20145 4385
rect 19829 4320 19835 4384
rect 19899 4320 19915 4384
rect 19979 4320 19995 4384
rect 20059 4320 20075 4384
rect 20139 4320 20145 4384
rect 19829 4319 20145 4320
rect 27603 4384 27919 4385
rect 27603 4320 27609 4384
rect 27673 4320 27689 4384
rect 27753 4320 27769 4384
rect 27833 4320 27849 4384
rect 27913 4320 27919 4384
rect 27603 4319 27919 4320
rect 8168 3840 8484 3841
rect 8168 3776 8174 3840
rect 8238 3776 8254 3840
rect 8318 3776 8334 3840
rect 8398 3776 8414 3840
rect 8478 3776 8484 3840
rect 8168 3775 8484 3776
rect 15942 3840 16258 3841
rect 15942 3776 15948 3840
rect 16012 3776 16028 3840
rect 16092 3776 16108 3840
rect 16172 3776 16188 3840
rect 16252 3776 16258 3840
rect 15942 3775 16258 3776
rect 23716 3840 24032 3841
rect 23716 3776 23722 3840
rect 23786 3776 23802 3840
rect 23866 3776 23882 3840
rect 23946 3776 23962 3840
rect 24026 3776 24032 3840
rect 23716 3775 24032 3776
rect 31490 3840 31806 3841
rect 31490 3776 31496 3840
rect 31560 3776 31576 3840
rect 31640 3776 31656 3840
rect 31720 3776 31736 3840
rect 31800 3776 31806 3840
rect 31490 3775 31806 3776
rect 4281 3296 4597 3297
rect 4281 3232 4287 3296
rect 4351 3232 4367 3296
rect 4431 3232 4447 3296
rect 4511 3232 4527 3296
rect 4591 3232 4597 3296
rect 4281 3231 4597 3232
rect 12055 3296 12371 3297
rect 12055 3232 12061 3296
rect 12125 3232 12141 3296
rect 12205 3232 12221 3296
rect 12285 3232 12301 3296
rect 12365 3232 12371 3296
rect 12055 3231 12371 3232
rect 19829 3296 20145 3297
rect 19829 3232 19835 3296
rect 19899 3232 19915 3296
rect 19979 3232 19995 3296
rect 20059 3232 20075 3296
rect 20139 3232 20145 3296
rect 19829 3231 20145 3232
rect 27603 3296 27919 3297
rect 27603 3232 27609 3296
rect 27673 3232 27689 3296
rect 27753 3232 27769 3296
rect 27833 3232 27849 3296
rect 27913 3232 27919 3296
rect 27603 3231 27919 3232
rect 8168 2752 8484 2753
rect 8168 2688 8174 2752
rect 8238 2688 8254 2752
rect 8318 2688 8334 2752
rect 8398 2688 8414 2752
rect 8478 2688 8484 2752
rect 8168 2687 8484 2688
rect 15942 2752 16258 2753
rect 15942 2688 15948 2752
rect 16012 2688 16028 2752
rect 16092 2688 16108 2752
rect 16172 2688 16188 2752
rect 16252 2688 16258 2752
rect 15942 2687 16258 2688
rect 23716 2752 24032 2753
rect 23716 2688 23722 2752
rect 23786 2688 23802 2752
rect 23866 2688 23882 2752
rect 23946 2688 23962 2752
rect 24026 2688 24032 2752
rect 23716 2687 24032 2688
rect 31490 2752 31806 2753
rect 31490 2688 31496 2752
rect 31560 2688 31576 2752
rect 31640 2688 31656 2752
rect 31720 2688 31736 2752
rect 31800 2688 31806 2752
rect 31490 2687 31806 2688
rect 4281 2208 4597 2209
rect 4281 2144 4287 2208
rect 4351 2144 4367 2208
rect 4431 2144 4447 2208
rect 4511 2144 4527 2208
rect 4591 2144 4597 2208
rect 4281 2143 4597 2144
rect 12055 2208 12371 2209
rect 12055 2144 12061 2208
rect 12125 2144 12141 2208
rect 12205 2144 12221 2208
rect 12285 2144 12301 2208
rect 12365 2144 12371 2208
rect 12055 2143 12371 2144
rect 19829 2208 20145 2209
rect 19829 2144 19835 2208
rect 19899 2144 19915 2208
rect 19979 2144 19995 2208
rect 20059 2144 20075 2208
rect 20139 2144 20145 2208
rect 19829 2143 20145 2144
rect 27603 2208 27919 2209
rect 27603 2144 27609 2208
rect 27673 2144 27689 2208
rect 27753 2144 27769 2208
rect 27833 2144 27849 2208
rect 27913 2144 27919 2208
rect 27603 2143 27919 2144
rect 8168 1664 8484 1665
rect 8168 1600 8174 1664
rect 8238 1600 8254 1664
rect 8318 1600 8334 1664
rect 8398 1600 8414 1664
rect 8478 1600 8484 1664
rect 8168 1599 8484 1600
rect 15942 1664 16258 1665
rect 15942 1600 15948 1664
rect 16012 1600 16028 1664
rect 16092 1600 16108 1664
rect 16172 1600 16188 1664
rect 16252 1600 16258 1664
rect 15942 1599 16258 1600
rect 23716 1664 24032 1665
rect 23716 1600 23722 1664
rect 23786 1600 23802 1664
rect 23866 1600 23882 1664
rect 23946 1600 23962 1664
rect 24026 1600 24032 1664
rect 23716 1599 24032 1600
rect 31490 1664 31806 1665
rect 31490 1600 31496 1664
rect 31560 1600 31576 1664
rect 31640 1600 31656 1664
rect 31720 1600 31736 1664
rect 31800 1600 31806 1664
rect 31490 1599 31806 1600
rect 4281 1120 4597 1121
rect 4281 1056 4287 1120
rect 4351 1056 4367 1120
rect 4431 1056 4447 1120
rect 4511 1056 4527 1120
rect 4591 1056 4597 1120
rect 4281 1055 4597 1056
rect 12055 1120 12371 1121
rect 12055 1056 12061 1120
rect 12125 1056 12141 1120
rect 12205 1056 12221 1120
rect 12285 1056 12301 1120
rect 12365 1056 12371 1120
rect 12055 1055 12371 1056
rect 19829 1120 20145 1121
rect 19829 1056 19835 1120
rect 19899 1056 19915 1120
rect 19979 1056 19995 1120
rect 20059 1056 20075 1120
rect 20139 1056 20145 1120
rect 19829 1055 20145 1056
rect 27603 1120 27919 1121
rect 27603 1056 27609 1120
rect 27673 1056 27689 1120
rect 27753 1056 27769 1120
rect 27833 1056 27849 1120
rect 27913 1056 27919 1120
rect 27603 1055 27919 1056
rect 8168 576 8484 577
rect 8168 512 8174 576
rect 8238 512 8254 576
rect 8318 512 8334 576
rect 8398 512 8414 576
rect 8478 512 8484 576
rect 8168 511 8484 512
rect 15942 576 16258 577
rect 15942 512 15948 576
rect 16012 512 16028 576
rect 16092 512 16108 576
rect 16172 512 16188 576
rect 16252 512 16258 576
rect 15942 511 16258 512
rect 23716 576 24032 577
rect 23716 512 23722 576
rect 23786 512 23802 576
rect 23866 512 23882 576
rect 23946 512 23962 576
rect 24026 512 24032 576
rect 23716 511 24032 512
rect 31490 576 31806 577
rect 31490 512 31496 576
rect 31560 512 31576 576
rect 31640 512 31656 576
rect 31720 512 31736 576
rect 31800 512 31806 576
rect 31490 511 31806 512
<< via3 >>
rect 28948 22204 29012 22268
rect 4476 21992 4540 21996
rect 4476 21936 4526 21992
rect 4526 21936 4540 21992
rect 4476 21932 4540 21936
rect 8156 21932 8220 21996
rect 16252 21992 16316 21996
rect 16252 21936 16302 21992
rect 16302 21936 16316 21992
rect 16252 21932 16316 21936
rect 796 21856 860 21860
rect 796 21800 846 21856
rect 846 21800 860 21856
rect 796 21796 860 21800
rect 1532 21856 1596 21860
rect 1532 21800 1582 21856
rect 1582 21800 1596 21856
rect 1532 21796 1596 21800
rect 2268 21856 2332 21860
rect 2268 21800 2318 21856
rect 2318 21800 2332 21856
rect 2268 21796 2332 21800
rect 3004 21796 3068 21860
rect 3740 21856 3804 21860
rect 3740 21800 3790 21856
rect 3790 21800 3804 21856
rect 3740 21796 3804 21800
rect 5212 21856 5276 21860
rect 5212 21800 5262 21856
rect 5262 21800 5276 21856
rect 5212 21796 5276 21800
rect 5948 21856 6012 21860
rect 5948 21800 5998 21856
rect 5998 21800 6012 21856
rect 5948 21796 6012 21800
rect 6684 21856 6748 21860
rect 6684 21800 6734 21856
rect 6734 21800 6748 21856
rect 6684 21796 6748 21800
rect 7420 21856 7484 21860
rect 7420 21800 7470 21856
rect 7470 21800 7484 21856
rect 7420 21796 7484 21800
rect 8892 21856 8956 21860
rect 8892 21800 8942 21856
rect 8942 21800 8956 21856
rect 8892 21796 8956 21800
rect 9628 21856 9692 21860
rect 9628 21800 9678 21856
rect 9678 21800 9692 21856
rect 9628 21796 9692 21800
rect 10364 21856 10428 21860
rect 10364 21800 10414 21856
rect 10414 21800 10428 21856
rect 10364 21796 10428 21800
rect 11100 21856 11164 21860
rect 11100 21800 11150 21856
rect 11150 21800 11164 21856
rect 11100 21796 11164 21800
rect 11836 21856 11900 21860
rect 11836 21800 11886 21856
rect 11886 21800 11900 21856
rect 11836 21796 11900 21800
rect 12572 21856 12636 21860
rect 12572 21800 12622 21856
rect 12622 21800 12636 21856
rect 12572 21796 12636 21800
rect 13308 21796 13372 21860
rect 14044 21856 14108 21860
rect 14044 21800 14094 21856
rect 14094 21800 14108 21856
rect 14044 21796 14108 21800
rect 14780 21856 14844 21860
rect 14780 21800 14830 21856
rect 14830 21800 14844 21856
rect 14780 21796 14844 21800
rect 15516 21856 15580 21860
rect 15516 21800 15566 21856
rect 15566 21800 15580 21856
rect 15516 21796 15580 21800
rect 16988 21856 17052 21860
rect 16988 21800 17038 21856
rect 17038 21800 17052 21856
rect 16988 21796 17052 21800
rect 29500 21796 29564 21860
rect 4287 21788 4351 21792
rect 4287 21732 4291 21788
rect 4291 21732 4347 21788
rect 4347 21732 4351 21788
rect 4287 21728 4351 21732
rect 4367 21788 4431 21792
rect 4367 21732 4371 21788
rect 4371 21732 4427 21788
rect 4427 21732 4431 21788
rect 4367 21728 4431 21732
rect 4447 21788 4511 21792
rect 4447 21732 4451 21788
rect 4451 21732 4507 21788
rect 4507 21732 4511 21788
rect 4447 21728 4511 21732
rect 4527 21788 4591 21792
rect 4527 21732 4531 21788
rect 4531 21732 4587 21788
rect 4587 21732 4591 21788
rect 4527 21728 4591 21732
rect 12061 21788 12125 21792
rect 12061 21732 12065 21788
rect 12065 21732 12121 21788
rect 12121 21732 12125 21788
rect 12061 21728 12125 21732
rect 12141 21788 12205 21792
rect 12141 21732 12145 21788
rect 12145 21732 12201 21788
rect 12201 21732 12205 21788
rect 12141 21728 12205 21732
rect 12221 21788 12285 21792
rect 12221 21732 12225 21788
rect 12225 21732 12281 21788
rect 12281 21732 12285 21788
rect 12221 21728 12285 21732
rect 12301 21788 12365 21792
rect 12301 21732 12305 21788
rect 12305 21732 12361 21788
rect 12361 21732 12365 21788
rect 12301 21728 12365 21732
rect 19835 21788 19899 21792
rect 19835 21732 19839 21788
rect 19839 21732 19895 21788
rect 19895 21732 19899 21788
rect 19835 21728 19899 21732
rect 19915 21788 19979 21792
rect 19915 21732 19919 21788
rect 19919 21732 19975 21788
rect 19975 21732 19979 21788
rect 19915 21728 19979 21732
rect 19995 21788 20059 21792
rect 19995 21732 19999 21788
rect 19999 21732 20055 21788
rect 20055 21732 20059 21788
rect 19995 21728 20059 21732
rect 20075 21788 20139 21792
rect 20075 21732 20079 21788
rect 20079 21732 20135 21788
rect 20135 21732 20139 21788
rect 20075 21728 20139 21732
rect 27609 21788 27673 21792
rect 27609 21732 27613 21788
rect 27613 21732 27669 21788
rect 27669 21732 27673 21788
rect 27609 21728 27673 21732
rect 27689 21788 27753 21792
rect 27689 21732 27693 21788
rect 27693 21732 27749 21788
rect 27749 21732 27753 21788
rect 27689 21728 27753 21732
rect 27769 21788 27833 21792
rect 27769 21732 27773 21788
rect 27773 21732 27829 21788
rect 27829 21732 27833 21788
rect 27769 21728 27833 21732
rect 27849 21788 27913 21792
rect 27849 21732 27853 21788
rect 27853 21732 27909 21788
rect 27909 21732 27913 21788
rect 27849 21728 27913 21732
rect 8174 21244 8238 21248
rect 8174 21188 8178 21244
rect 8178 21188 8234 21244
rect 8234 21188 8238 21244
rect 8174 21184 8238 21188
rect 8254 21244 8318 21248
rect 8254 21188 8258 21244
rect 8258 21188 8314 21244
rect 8314 21188 8318 21244
rect 8254 21184 8318 21188
rect 8334 21244 8398 21248
rect 8334 21188 8338 21244
rect 8338 21188 8394 21244
rect 8394 21188 8398 21244
rect 8334 21184 8398 21188
rect 8414 21244 8478 21248
rect 8414 21188 8418 21244
rect 8418 21188 8474 21244
rect 8474 21188 8478 21244
rect 8414 21184 8478 21188
rect 15948 21244 16012 21248
rect 15948 21188 15952 21244
rect 15952 21188 16008 21244
rect 16008 21188 16012 21244
rect 15948 21184 16012 21188
rect 16028 21244 16092 21248
rect 16028 21188 16032 21244
rect 16032 21188 16088 21244
rect 16088 21188 16092 21244
rect 16028 21184 16092 21188
rect 16108 21244 16172 21248
rect 16108 21188 16112 21244
rect 16112 21188 16168 21244
rect 16168 21188 16172 21244
rect 16108 21184 16172 21188
rect 16188 21244 16252 21248
rect 16188 21188 16192 21244
rect 16192 21188 16248 21244
rect 16248 21188 16252 21244
rect 16188 21184 16252 21188
rect 23722 21244 23786 21248
rect 23722 21188 23726 21244
rect 23726 21188 23782 21244
rect 23782 21188 23786 21244
rect 23722 21184 23786 21188
rect 23802 21244 23866 21248
rect 23802 21188 23806 21244
rect 23806 21188 23862 21244
rect 23862 21188 23866 21244
rect 23802 21184 23866 21188
rect 23882 21244 23946 21248
rect 23882 21188 23886 21244
rect 23886 21188 23942 21244
rect 23942 21188 23946 21244
rect 23882 21184 23946 21188
rect 23962 21244 24026 21248
rect 23962 21188 23966 21244
rect 23966 21188 24022 21244
rect 24022 21188 24026 21244
rect 23962 21184 24026 21188
rect 31496 21244 31560 21248
rect 31496 21188 31500 21244
rect 31500 21188 31556 21244
rect 31556 21188 31560 21244
rect 31496 21184 31560 21188
rect 31576 21244 31640 21248
rect 31576 21188 31580 21244
rect 31580 21188 31636 21244
rect 31636 21188 31640 21244
rect 31576 21184 31640 21188
rect 31656 21244 31720 21248
rect 31656 21188 31660 21244
rect 31660 21188 31716 21244
rect 31716 21188 31720 21244
rect 31656 21184 31720 21188
rect 31736 21244 31800 21248
rect 31736 21188 31740 21244
rect 31740 21188 31796 21244
rect 31796 21188 31800 21244
rect 31736 21184 31800 21188
rect 4287 20700 4351 20704
rect 4287 20644 4291 20700
rect 4291 20644 4347 20700
rect 4347 20644 4351 20700
rect 4287 20640 4351 20644
rect 4367 20700 4431 20704
rect 4367 20644 4371 20700
rect 4371 20644 4427 20700
rect 4427 20644 4431 20700
rect 4367 20640 4431 20644
rect 4447 20700 4511 20704
rect 4447 20644 4451 20700
rect 4451 20644 4507 20700
rect 4507 20644 4511 20700
rect 4447 20640 4511 20644
rect 4527 20700 4591 20704
rect 4527 20644 4531 20700
rect 4531 20644 4587 20700
rect 4587 20644 4591 20700
rect 4527 20640 4591 20644
rect 12061 20700 12125 20704
rect 12061 20644 12065 20700
rect 12065 20644 12121 20700
rect 12121 20644 12125 20700
rect 12061 20640 12125 20644
rect 12141 20700 12205 20704
rect 12141 20644 12145 20700
rect 12145 20644 12201 20700
rect 12201 20644 12205 20700
rect 12141 20640 12205 20644
rect 12221 20700 12285 20704
rect 12221 20644 12225 20700
rect 12225 20644 12281 20700
rect 12281 20644 12285 20700
rect 12221 20640 12285 20644
rect 12301 20700 12365 20704
rect 12301 20644 12305 20700
rect 12305 20644 12361 20700
rect 12361 20644 12365 20700
rect 12301 20640 12365 20644
rect 19835 20700 19899 20704
rect 19835 20644 19839 20700
rect 19839 20644 19895 20700
rect 19895 20644 19899 20700
rect 19835 20640 19899 20644
rect 19915 20700 19979 20704
rect 19915 20644 19919 20700
rect 19919 20644 19975 20700
rect 19975 20644 19979 20700
rect 19915 20640 19979 20644
rect 19995 20700 20059 20704
rect 19995 20644 19999 20700
rect 19999 20644 20055 20700
rect 20055 20644 20059 20700
rect 19995 20640 20059 20644
rect 20075 20700 20139 20704
rect 20075 20644 20079 20700
rect 20079 20644 20135 20700
rect 20135 20644 20139 20700
rect 20075 20640 20139 20644
rect 27609 20700 27673 20704
rect 27609 20644 27613 20700
rect 27613 20644 27669 20700
rect 27669 20644 27673 20700
rect 27609 20640 27673 20644
rect 27689 20700 27753 20704
rect 27689 20644 27693 20700
rect 27693 20644 27749 20700
rect 27749 20644 27753 20700
rect 27689 20640 27753 20644
rect 27769 20700 27833 20704
rect 27769 20644 27773 20700
rect 27773 20644 27829 20700
rect 27829 20644 27833 20700
rect 27769 20640 27833 20644
rect 27849 20700 27913 20704
rect 27849 20644 27853 20700
rect 27853 20644 27909 20700
rect 27909 20644 27913 20700
rect 27849 20640 27913 20644
rect 8174 20156 8238 20160
rect 8174 20100 8178 20156
rect 8178 20100 8234 20156
rect 8234 20100 8238 20156
rect 8174 20096 8238 20100
rect 8254 20156 8318 20160
rect 8254 20100 8258 20156
rect 8258 20100 8314 20156
rect 8314 20100 8318 20156
rect 8254 20096 8318 20100
rect 8334 20156 8398 20160
rect 8334 20100 8338 20156
rect 8338 20100 8394 20156
rect 8394 20100 8398 20156
rect 8334 20096 8398 20100
rect 8414 20156 8478 20160
rect 8414 20100 8418 20156
rect 8418 20100 8474 20156
rect 8474 20100 8478 20156
rect 8414 20096 8478 20100
rect 15948 20156 16012 20160
rect 15948 20100 15952 20156
rect 15952 20100 16008 20156
rect 16008 20100 16012 20156
rect 15948 20096 16012 20100
rect 16028 20156 16092 20160
rect 16028 20100 16032 20156
rect 16032 20100 16088 20156
rect 16088 20100 16092 20156
rect 16028 20096 16092 20100
rect 16108 20156 16172 20160
rect 16108 20100 16112 20156
rect 16112 20100 16168 20156
rect 16168 20100 16172 20156
rect 16108 20096 16172 20100
rect 16188 20156 16252 20160
rect 16188 20100 16192 20156
rect 16192 20100 16248 20156
rect 16248 20100 16252 20156
rect 16188 20096 16252 20100
rect 23722 20156 23786 20160
rect 23722 20100 23726 20156
rect 23726 20100 23782 20156
rect 23782 20100 23786 20156
rect 23722 20096 23786 20100
rect 23802 20156 23866 20160
rect 23802 20100 23806 20156
rect 23806 20100 23862 20156
rect 23862 20100 23866 20156
rect 23802 20096 23866 20100
rect 23882 20156 23946 20160
rect 23882 20100 23886 20156
rect 23886 20100 23942 20156
rect 23942 20100 23946 20156
rect 23882 20096 23946 20100
rect 23962 20156 24026 20160
rect 23962 20100 23966 20156
rect 23966 20100 24022 20156
rect 24022 20100 24026 20156
rect 23962 20096 24026 20100
rect 31496 20156 31560 20160
rect 31496 20100 31500 20156
rect 31500 20100 31556 20156
rect 31556 20100 31560 20156
rect 31496 20096 31560 20100
rect 31576 20156 31640 20160
rect 31576 20100 31580 20156
rect 31580 20100 31636 20156
rect 31636 20100 31640 20156
rect 31576 20096 31640 20100
rect 31656 20156 31720 20160
rect 31656 20100 31660 20156
rect 31660 20100 31716 20156
rect 31716 20100 31720 20156
rect 31656 20096 31720 20100
rect 31736 20156 31800 20160
rect 31736 20100 31740 20156
rect 31740 20100 31796 20156
rect 31796 20100 31800 20156
rect 31736 20096 31800 20100
rect 4287 19612 4351 19616
rect 4287 19556 4291 19612
rect 4291 19556 4347 19612
rect 4347 19556 4351 19612
rect 4287 19552 4351 19556
rect 4367 19612 4431 19616
rect 4367 19556 4371 19612
rect 4371 19556 4427 19612
rect 4427 19556 4431 19612
rect 4367 19552 4431 19556
rect 4447 19612 4511 19616
rect 4447 19556 4451 19612
rect 4451 19556 4507 19612
rect 4507 19556 4511 19612
rect 4447 19552 4511 19556
rect 4527 19612 4591 19616
rect 4527 19556 4531 19612
rect 4531 19556 4587 19612
rect 4587 19556 4591 19612
rect 4527 19552 4591 19556
rect 12061 19612 12125 19616
rect 12061 19556 12065 19612
rect 12065 19556 12121 19612
rect 12121 19556 12125 19612
rect 12061 19552 12125 19556
rect 12141 19612 12205 19616
rect 12141 19556 12145 19612
rect 12145 19556 12201 19612
rect 12201 19556 12205 19612
rect 12141 19552 12205 19556
rect 12221 19612 12285 19616
rect 12221 19556 12225 19612
rect 12225 19556 12281 19612
rect 12281 19556 12285 19612
rect 12221 19552 12285 19556
rect 12301 19612 12365 19616
rect 12301 19556 12305 19612
rect 12305 19556 12361 19612
rect 12361 19556 12365 19612
rect 12301 19552 12365 19556
rect 19835 19612 19899 19616
rect 19835 19556 19839 19612
rect 19839 19556 19895 19612
rect 19895 19556 19899 19612
rect 19835 19552 19899 19556
rect 19915 19612 19979 19616
rect 19915 19556 19919 19612
rect 19919 19556 19975 19612
rect 19975 19556 19979 19612
rect 19915 19552 19979 19556
rect 19995 19612 20059 19616
rect 19995 19556 19999 19612
rect 19999 19556 20055 19612
rect 20055 19556 20059 19612
rect 19995 19552 20059 19556
rect 20075 19612 20139 19616
rect 20075 19556 20079 19612
rect 20079 19556 20135 19612
rect 20135 19556 20139 19612
rect 20075 19552 20139 19556
rect 27609 19612 27673 19616
rect 27609 19556 27613 19612
rect 27613 19556 27669 19612
rect 27669 19556 27673 19612
rect 27609 19552 27673 19556
rect 27689 19612 27753 19616
rect 27689 19556 27693 19612
rect 27693 19556 27749 19612
rect 27749 19556 27753 19612
rect 27689 19552 27753 19556
rect 27769 19612 27833 19616
rect 27769 19556 27773 19612
rect 27773 19556 27829 19612
rect 27829 19556 27833 19612
rect 27769 19552 27833 19556
rect 27849 19612 27913 19616
rect 27849 19556 27853 19612
rect 27853 19556 27909 19612
rect 27909 19556 27913 19612
rect 27849 19552 27913 19556
rect 17724 19212 17788 19276
rect 8174 19068 8238 19072
rect 8174 19012 8178 19068
rect 8178 19012 8234 19068
rect 8234 19012 8238 19068
rect 8174 19008 8238 19012
rect 8254 19068 8318 19072
rect 8254 19012 8258 19068
rect 8258 19012 8314 19068
rect 8314 19012 8318 19068
rect 8254 19008 8318 19012
rect 8334 19068 8398 19072
rect 8334 19012 8338 19068
rect 8338 19012 8394 19068
rect 8394 19012 8398 19068
rect 8334 19008 8398 19012
rect 8414 19068 8478 19072
rect 8414 19012 8418 19068
rect 8418 19012 8474 19068
rect 8474 19012 8478 19068
rect 8414 19008 8478 19012
rect 15948 19068 16012 19072
rect 15948 19012 15952 19068
rect 15952 19012 16008 19068
rect 16008 19012 16012 19068
rect 15948 19008 16012 19012
rect 16028 19068 16092 19072
rect 16028 19012 16032 19068
rect 16032 19012 16088 19068
rect 16088 19012 16092 19068
rect 16028 19008 16092 19012
rect 16108 19068 16172 19072
rect 16108 19012 16112 19068
rect 16112 19012 16168 19068
rect 16168 19012 16172 19068
rect 16108 19008 16172 19012
rect 16188 19068 16252 19072
rect 16188 19012 16192 19068
rect 16192 19012 16248 19068
rect 16248 19012 16252 19068
rect 16188 19008 16252 19012
rect 23722 19068 23786 19072
rect 23722 19012 23726 19068
rect 23726 19012 23782 19068
rect 23782 19012 23786 19068
rect 23722 19008 23786 19012
rect 23802 19068 23866 19072
rect 23802 19012 23806 19068
rect 23806 19012 23862 19068
rect 23862 19012 23866 19068
rect 23802 19008 23866 19012
rect 23882 19068 23946 19072
rect 23882 19012 23886 19068
rect 23886 19012 23942 19068
rect 23942 19012 23946 19068
rect 23882 19008 23946 19012
rect 23962 19068 24026 19072
rect 23962 19012 23966 19068
rect 23966 19012 24022 19068
rect 24022 19012 24026 19068
rect 23962 19008 24026 19012
rect 31496 19068 31560 19072
rect 31496 19012 31500 19068
rect 31500 19012 31556 19068
rect 31556 19012 31560 19068
rect 31496 19008 31560 19012
rect 31576 19068 31640 19072
rect 31576 19012 31580 19068
rect 31580 19012 31636 19068
rect 31636 19012 31640 19068
rect 31576 19008 31640 19012
rect 31656 19068 31720 19072
rect 31656 19012 31660 19068
rect 31660 19012 31716 19068
rect 31716 19012 31720 19068
rect 31656 19008 31720 19012
rect 31736 19068 31800 19072
rect 31736 19012 31740 19068
rect 31740 19012 31796 19068
rect 31796 19012 31800 19068
rect 31736 19008 31800 19012
rect 4287 18524 4351 18528
rect 4287 18468 4291 18524
rect 4291 18468 4347 18524
rect 4347 18468 4351 18524
rect 4287 18464 4351 18468
rect 4367 18524 4431 18528
rect 4367 18468 4371 18524
rect 4371 18468 4427 18524
rect 4427 18468 4431 18524
rect 4367 18464 4431 18468
rect 4447 18524 4511 18528
rect 4447 18468 4451 18524
rect 4451 18468 4507 18524
rect 4507 18468 4511 18524
rect 4447 18464 4511 18468
rect 4527 18524 4591 18528
rect 4527 18468 4531 18524
rect 4531 18468 4587 18524
rect 4587 18468 4591 18524
rect 4527 18464 4591 18468
rect 12061 18524 12125 18528
rect 12061 18468 12065 18524
rect 12065 18468 12121 18524
rect 12121 18468 12125 18524
rect 12061 18464 12125 18468
rect 12141 18524 12205 18528
rect 12141 18468 12145 18524
rect 12145 18468 12201 18524
rect 12201 18468 12205 18524
rect 12141 18464 12205 18468
rect 12221 18524 12285 18528
rect 12221 18468 12225 18524
rect 12225 18468 12281 18524
rect 12281 18468 12285 18524
rect 12221 18464 12285 18468
rect 12301 18524 12365 18528
rect 12301 18468 12305 18524
rect 12305 18468 12361 18524
rect 12361 18468 12365 18524
rect 12301 18464 12365 18468
rect 19835 18524 19899 18528
rect 19835 18468 19839 18524
rect 19839 18468 19895 18524
rect 19895 18468 19899 18524
rect 19835 18464 19899 18468
rect 19915 18524 19979 18528
rect 19915 18468 19919 18524
rect 19919 18468 19975 18524
rect 19975 18468 19979 18524
rect 19915 18464 19979 18468
rect 19995 18524 20059 18528
rect 19995 18468 19999 18524
rect 19999 18468 20055 18524
rect 20055 18468 20059 18524
rect 19995 18464 20059 18468
rect 20075 18524 20139 18528
rect 20075 18468 20079 18524
rect 20079 18468 20135 18524
rect 20135 18468 20139 18524
rect 20075 18464 20139 18468
rect 27609 18524 27673 18528
rect 27609 18468 27613 18524
rect 27613 18468 27669 18524
rect 27669 18468 27673 18524
rect 27609 18464 27673 18468
rect 27689 18524 27753 18528
rect 27689 18468 27693 18524
rect 27693 18468 27749 18524
rect 27749 18468 27753 18524
rect 27689 18464 27753 18468
rect 27769 18524 27833 18528
rect 27769 18468 27773 18524
rect 27773 18468 27829 18524
rect 27829 18468 27833 18524
rect 27769 18464 27833 18468
rect 27849 18524 27913 18528
rect 27849 18468 27853 18524
rect 27853 18468 27909 18524
rect 27909 18468 27913 18524
rect 27849 18464 27913 18468
rect 8174 17980 8238 17984
rect 8174 17924 8178 17980
rect 8178 17924 8234 17980
rect 8234 17924 8238 17980
rect 8174 17920 8238 17924
rect 8254 17980 8318 17984
rect 8254 17924 8258 17980
rect 8258 17924 8314 17980
rect 8314 17924 8318 17980
rect 8254 17920 8318 17924
rect 8334 17980 8398 17984
rect 8334 17924 8338 17980
rect 8338 17924 8394 17980
rect 8394 17924 8398 17980
rect 8334 17920 8398 17924
rect 8414 17980 8478 17984
rect 8414 17924 8418 17980
rect 8418 17924 8474 17980
rect 8474 17924 8478 17980
rect 8414 17920 8478 17924
rect 15948 17980 16012 17984
rect 15948 17924 15952 17980
rect 15952 17924 16008 17980
rect 16008 17924 16012 17980
rect 15948 17920 16012 17924
rect 16028 17980 16092 17984
rect 16028 17924 16032 17980
rect 16032 17924 16088 17980
rect 16088 17924 16092 17980
rect 16028 17920 16092 17924
rect 16108 17980 16172 17984
rect 16108 17924 16112 17980
rect 16112 17924 16168 17980
rect 16168 17924 16172 17980
rect 16108 17920 16172 17924
rect 16188 17980 16252 17984
rect 16188 17924 16192 17980
rect 16192 17924 16248 17980
rect 16248 17924 16252 17980
rect 16188 17920 16252 17924
rect 23722 17980 23786 17984
rect 23722 17924 23726 17980
rect 23726 17924 23782 17980
rect 23782 17924 23786 17980
rect 23722 17920 23786 17924
rect 23802 17980 23866 17984
rect 23802 17924 23806 17980
rect 23806 17924 23862 17980
rect 23862 17924 23866 17980
rect 23802 17920 23866 17924
rect 23882 17980 23946 17984
rect 23882 17924 23886 17980
rect 23886 17924 23942 17980
rect 23942 17924 23946 17980
rect 23882 17920 23946 17924
rect 23962 17980 24026 17984
rect 23962 17924 23966 17980
rect 23966 17924 24022 17980
rect 24022 17924 24026 17980
rect 23962 17920 24026 17924
rect 31496 17980 31560 17984
rect 31496 17924 31500 17980
rect 31500 17924 31556 17980
rect 31556 17924 31560 17980
rect 31496 17920 31560 17924
rect 31576 17980 31640 17984
rect 31576 17924 31580 17980
rect 31580 17924 31636 17980
rect 31636 17924 31640 17980
rect 31576 17920 31640 17924
rect 31656 17980 31720 17984
rect 31656 17924 31660 17980
rect 31660 17924 31716 17980
rect 31716 17924 31720 17980
rect 31656 17920 31720 17924
rect 31736 17980 31800 17984
rect 31736 17924 31740 17980
rect 31740 17924 31796 17980
rect 31796 17924 31800 17980
rect 31736 17920 31800 17924
rect 4287 17436 4351 17440
rect 4287 17380 4291 17436
rect 4291 17380 4347 17436
rect 4347 17380 4351 17436
rect 4287 17376 4351 17380
rect 4367 17436 4431 17440
rect 4367 17380 4371 17436
rect 4371 17380 4427 17436
rect 4427 17380 4431 17436
rect 4367 17376 4431 17380
rect 4447 17436 4511 17440
rect 4447 17380 4451 17436
rect 4451 17380 4507 17436
rect 4507 17380 4511 17436
rect 4447 17376 4511 17380
rect 4527 17436 4591 17440
rect 4527 17380 4531 17436
rect 4531 17380 4587 17436
rect 4587 17380 4591 17436
rect 4527 17376 4591 17380
rect 12061 17436 12125 17440
rect 12061 17380 12065 17436
rect 12065 17380 12121 17436
rect 12121 17380 12125 17436
rect 12061 17376 12125 17380
rect 12141 17436 12205 17440
rect 12141 17380 12145 17436
rect 12145 17380 12201 17436
rect 12201 17380 12205 17436
rect 12141 17376 12205 17380
rect 12221 17436 12285 17440
rect 12221 17380 12225 17436
rect 12225 17380 12281 17436
rect 12281 17380 12285 17436
rect 12221 17376 12285 17380
rect 12301 17436 12365 17440
rect 12301 17380 12305 17436
rect 12305 17380 12361 17436
rect 12361 17380 12365 17436
rect 12301 17376 12365 17380
rect 19835 17436 19899 17440
rect 19835 17380 19839 17436
rect 19839 17380 19895 17436
rect 19895 17380 19899 17436
rect 19835 17376 19899 17380
rect 19915 17436 19979 17440
rect 19915 17380 19919 17436
rect 19919 17380 19975 17436
rect 19975 17380 19979 17436
rect 19915 17376 19979 17380
rect 19995 17436 20059 17440
rect 19995 17380 19999 17436
rect 19999 17380 20055 17436
rect 20055 17380 20059 17436
rect 19995 17376 20059 17380
rect 20075 17436 20139 17440
rect 20075 17380 20079 17436
rect 20079 17380 20135 17436
rect 20135 17380 20139 17436
rect 20075 17376 20139 17380
rect 27609 17436 27673 17440
rect 27609 17380 27613 17436
rect 27613 17380 27669 17436
rect 27669 17380 27673 17436
rect 27609 17376 27673 17380
rect 27689 17436 27753 17440
rect 27689 17380 27693 17436
rect 27693 17380 27749 17436
rect 27749 17380 27753 17436
rect 27689 17376 27753 17380
rect 27769 17436 27833 17440
rect 27769 17380 27773 17436
rect 27773 17380 27829 17436
rect 27829 17380 27833 17436
rect 27769 17376 27833 17380
rect 27849 17436 27913 17440
rect 27849 17380 27853 17436
rect 27853 17380 27909 17436
rect 27909 17380 27913 17436
rect 27849 17376 27913 17380
rect 8174 16892 8238 16896
rect 8174 16836 8178 16892
rect 8178 16836 8234 16892
rect 8234 16836 8238 16892
rect 8174 16832 8238 16836
rect 8254 16892 8318 16896
rect 8254 16836 8258 16892
rect 8258 16836 8314 16892
rect 8314 16836 8318 16892
rect 8254 16832 8318 16836
rect 8334 16892 8398 16896
rect 8334 16836 8338 16892
rect 8338 16836 8394 16892
rect 8394 16836 8398 16892
rect 8334 16832 8398 16836
rect 8414 16892 8478 16896
rect 8414 16836 8418 16892
rect 8418 16836 8474 16892
rect 8474 16836 8478 16892
rect 8414 16832 8478 16836
rect 15948 16892 16012 16896
rect 15948 16836 15952 16892
rect 15952 16836 16008 16892
rect 16008 16836 16012 16892
rect 15948 16832 16012 16836
rect 16028 16892 16092 16896
rect 16028 16836 16032 16892
rect 16032 16836 16088 16892
rect 16088 16836 16092 16892
rect 16028 16832 16092 16836
rect 16108 16892 16172 16896
rect 16108 16836 16112 16892
rect 16112 16836 16168 16892
rect 16168 16836 16172 16892
rect 16108 16832 16172 16836
rect 16188 16892 16252 16896
rect 16188 16836 16192 16892
rect 16192 16836 16248 16892
rect 16248 16836 16252 16892
rect 16188 16832 16252 16836
rect 23722 16892 23786 16896
rect 23722 16836 23726 16892
rect 23726 16836 23782 16892
rect 23782 16836 23786 16892
rect 23722 16832 23786 16836
rect 23802 16892 23866 16896
rect 23802 16836 23806 16892
rect 23806 16836 23862 16892
rect 23862 16836 23866 16892
rect 23802 16832 23866 16836
rect 23882 16892 23946 16896
rect 23882 16836 23886 16892
rect 23886 16836 23942 16892
rect 23942 16836 23946 16892
rect 23882 16832 23946 16836
rect 23962 16892 24026 16896
rect 23962 16836 23966 16892
rect 23966 16836 24022 16892
rect 24022 16836 24026 16892
rect 23962 16832 24026 16836
rect 31496 16892 31560 16896
rect 31496 16836 31500 16892
rect 31500 16836 31556 16892
rect 31556 16836 31560 16892
rect 31496 16832 31560 16836
rect 31576 16892 31640 16896
rect 31576 16836 31580 16892
rect 31580 16836 31636 16892
rect 31636 16836 31640 16892
rect 31576 16832 31640 16836
rect 31656 16892 31720 16896
rect 31656 16836 31660 16892
rect 31660 16836 31716 16892
rect 31716 16836 31720 16892
rect 31656 16832 31720 16836
rect 31736 16892 31800 16896
rect 31736 16836 31740 16892
rect 31740 16836 31796 16892
rect 31796 16836 31800 16892
rect 31736 16832 31800 16836
rect 4287 16348 4351 16352
rect 4287 16292 4291 16348
rect 4291 16292 4347 16348
rect 4347 16292 4351 16348
rect 4287 16288 4351 16292
rect 4367 16348 4431 16352
rect 4367 16292 4371 16348
rect 4371 16292 4427 16348
rect 4427 16292 4431 16348
rect 4367 16288 4431 16292
rect 4447 16348 4511 16352
rect 4447 16292 4451 16348
rect 4451 16292 4507 16348
rect 4507 16292 4511 16348
rect 4447 16288 4511 16292
rect 4527 16348 4591 16352
rect 4527 16292 4531 16348
rect 4531 16292 4587 16348
rect 4587 16292 4591 16348
rect 4527 16288 4591 16292
rect 12061 16348 12125 16352
rect 12061 16292 12065 16348
rect 12065 16292 12121 16348
rect 12121 16292 12125 16348
rect 12061 16288 12125 16292
rect 12141 16348 12205 16352
rect 12141 16292 12145 16348
rect 12145 16292 12201 16348
rect 12201 16292 12205 16348
rect 12141 16288 12205 16292
rect 12221 16348 12285 16352
rect 12221 16292 12225 16348
rect 12225 16292 12281 16348
rect 12281 16292 12285 16348
rect 12221 16288 12285 16292
rect 12301 16348 12365 16352
rect 12301 16292 12305 16348
rect 12305 16292 12361 16348
rect 12361 16292 12365 16348
rect 12301 16288 12365 16292
rect 19835 16348 19899 16352
rect 19835 16292 19839 16348
rect 19839 16292 19895 16348
rect 19895 16292 19899 16348
rect 19835 16288 19899 16292
rect 19915 16348 19979 16352
rect 19915 16292 19919 16348
rect 19919 16292 19975 16348
rect 19975 16292 19979 16348
rect 19915 16288 19979 16292
rect 19995 16348 20059 16352
rect 19995 16292 19999 16348
rect 19999 16292 20055 16348
rect 20055 16292 20059 16348
rect 19995 16288 20059 16292
rect 20075 16348 20139 16352
rect 20075 16292 20079 16348
rect 20079 16292 20135 16348
rect 20135 16292 20139 16348
rect 20075 16288 20139 16292
rect 27609 16348 27673 16352
rect 27609 16292 27613 16348
rect 27613 16292 27669 16348
rect 27669 16292 27673 16348
rect 27609 16288 27673 16292
rect 27689 16348 27753 16352
rect 27689 16292 27693 16348
rect 27693 16292 27749 16348
rect 27749 16292 27753 16348
rect 27689 16288 27753 16292
rect 27769 16348 27833 16352
rect 27769 16292 27773 16348
rect 27773 16292 27829 16348
rect 27829 16292 27833 16348
rect 27769 16288 27833 16292
rect 27849 16348 27913 16352
rect 27849 16292 27853 16348
rect 27853 16292 27909 16348
rect 27909 16292 27913 16348
rect 27849 16288 27913 16292
rect 8174 15804 8238 15808
rect 8174 15748 8178 15804
rect 8178 15748 8234 15804
rect 8234 15748 8238 15804
rect 8174 15744 8238 15748
rect 8254 15804 8318 15808
rect 8254 15748 8258 15804
rect 8258 15748 8314 15804
rect 8314 15748 8318 15804
rect 8254 15744 8318 15748
rect 8334 15804 8398 15808
rect 8334 15748 8338 15804
rect 8338 15748 8394 15804
rect 8394 15748 8398 15804
rect 8334 15744 8398 15748
rect 8414 15804 8478 15808
rect 8414 15748 8418 15804
rect 8418 15748 8474 15804
rect 8474 15748 8478 15804
rect 8414 15744 8478 15748
rect 15948 15804 16012 15808
rect 15948 15748 15952 15804
rect 15952 15748 16008 15804
rect 16008 15748 16012 15804
rect 15948 15744 16012 15748
rect 16028 15804 16092 15808
rect 16028 15748 16032 15804
rect 16032 15748 16088 15804
rect 16088 15748 16092 15804
rect 16028 15744 16092 15748
rect 16108 15804 16172 15808
rect 16108 15748 16112 15804
rect 16112 15748 16168 15804
rect 16168 15748 16172 15804
rect 16108 15744 16172 15748
rect 16188 15804 16252 15808
rect 16188 15748 16192 15804
rect 16192 15748 16248 15804
rect 16248 15748 16252 15804
rect 16188 15744 16252 15748
rect 23722 15804 23786 15808
rect 23722 15748 23726 15804
rect 23726 15748 23782 15804
rect 23782 15748 23786 15804
rect 23722 15744 23786 15748
rect 23802 15804 23866 15808
rect 23802 15748 23806 15804
rect 23806 15748 23862 15804
rect 23862 15748 23866 15804
rect 23802 15744 23866 15748
rect 23882 15804 23946 15808
rect 23882 15748 23886 15804
rect 23886 15748 23942 15804
rect 23942 15748 23946 15804
rect 23882 15744 23946 15748
rect 23962 15804 24026 15808
rect 23962 15748 23966 15804
rect 23966 15748 24022 15804
rect 24022 15748 24026 15804
rect 23962 15744 24026 15748
rect 31496 15804 31560 15808
rect 31496 15748 31500 15804
rect 31500 15748 31556 15804
rect 31556 15748 31560 15804
rect 31496 15744 31560 15748
rect 31576 15804 31640 15808
rect 31576 15748 31580 15804
rect 31580 15748 31636 15804
rect 31636 15748 31640 15804
rect 31576 15744 31640 15748
rect 31656 15804 31720 15808
rect 31656 15748 31660 15804
rect 31660 15748 31716 15804
rect 31716 15748 31720 15804
rect 31656 15744 31720 15748
rect 31736 15804 31800 15808
rect 31736 15748 31740 15804
rect 31740 15748 31796 15804
rect 31796 15748 31800 15804
rect 31736 15744 31800 15748
rect 4287 15260 4351 15264
rect 4287 15204 4291 15260
rect 4291 15204 4347 15260
rect 4347 15204 4351 15260
rect 4287 15200 4351 15204
rect 4367 15260 4431 15264
rect 4367 15204 4371 15260
rect 4371 15204 4427 15260
rect 4427 15204 4431 15260
rect 4367 15200 4431 15204
rect 4447 15260 4511 15264
rect 4447 15204 4451 15260
rect 4451 15204 4507 15260
rect 4507 15204 4511 15260
rect 4447 15200 4511 15204
rect 4527 15260 4591 15264
rect 4527 15204 4531 15260
rect 4531 15204 4587 15260
rect 4587 15204 4591 15260
rect 4527 15200 4591 15204
rect 12061 15260 12125 15264
rect 12061 15204 12065 15260
rect 12065 15204 12121 15260
rect 12121 15204 12125 15260
rect 12061 15200 12125 15204
rect 12141 15260 12205 15264
rect 12141 15204 12145 15260
rect 12145 15204 12201 15260
rect 12201 15204 12205 15260
rect 12141 15200 12205 15204
rect 12221 15260 12285 15264
rect 12221 15204 12225 15260
rect 12225 15204 12281 15260
rect 12281 15204 12285 15260
rect 12221 15200 12285 15204
rect 12301 15260 12365 15264
rect 12301 15204 12305 15260
rect 12305 15204 12361 15260
rect 12361 15204 12365 15260
rect 12301 15200 12365 15204
rect 19835 15260 19899 15264
rect 19835 15204 19839 15260
rect 19839 15204 19895 15260
rect 19895 15204 19899 15260
rect 19835 15200 19899 15204
rect 19915 15260 19979 15264
rect 19915 15204 19919 15260
rect 19919 15204 19975 15260
rect 19975 15204 19979 15260
rect 19915 15200 19979 15204
rect 19995 15260 20059 15264
rect 19995 15204 19999 15260
rect 19999 15204 20055 15260
rect 20055 15204 20059 15260
rect 19995 15200 20059 15204
rect 20075 15260 20139 15264
rect 20075 15204 20079 15260
rect 20079 15204 20135 15260
rect 20135 15204 20139 15260
rect 20075 15200 20139 15204
rect 27609 15260 27673 15264
rect 27609 15204 27613 15260
rect 27613 15204 27669 15260
rect 27669 15204 27673 15260
rect 27609 15200 27673 15204
rect 27689 15260 27753 15264
rect 27689 15204 27693 15260
rect 27693 15204 27749 15260
rect 27749 15204 27753 15260
rect 27689 15200 27753 15204
rect 27769 15260 27833 15264
rect 27769 15204 27773 15260
rect 27773 15204 27829 15260
rect 27829 15204 27833 15260
rect 27769 15200 27833 15204
rect 27849 15260 27913 15264
rect 27849 15204 27853 15260
rect 27853 15204 27909 15260
rect 27909 15204 27913 15260
rect 27849 15200 27913 15204
rect 8174 14716 8238 14720
rect 8174 14660 8178 14716
rect 8178 14660 8234 14716
rect 8234 14660 8238 14716
rect 8174 14656 8238 14660
rect 8254 14716 8318 14720
rect 8254 14660 8258 14716
rect 8258 14660 8314 14716
rect 8314 14660 8318 14716
rect 8254 14656 8318 14660
rect 8334 14716 8398 14720
rect 8334 14660 8338 14716
rect 8338 14660 8394 14716
rect 8394 14660 8398 14716
rect 8334 14656 8398 14660
rect 8414 14716 8478 14720
rect 8414 14660 8418 14716
rect 8418 14660 8474 14716
rect 8474 14660 8478 14716
rect 8414 14656 8478 14660
rect 15948 14716 16012 14720
rect 15948 14660 15952 14716
rect 15952 14660 16008 14716
rect 16008 14660 16012 14716
rect 15948 14656 16012 14660
rect 16028 14716 16092 14720
rect 16028 14660 16032 14716
rect 16032 14660 16088 14716
rect 16088 14660 16092 14716
rect 16028 14656 16092 14660
rect 16108 14716 16172 14720
rect 16108 14660 16112 14716
rect 16112 14660 16168 14716
rect 16168 14660 16172 14716
rect 16108 14656 16172 14660
rect 16188 14716 16252 14720
rect 16188 14660 16192 14716
rect 16192 14660 16248 14716
rect 16248 14660 16252 14716
rect 16188 14656 16252 14660
rect 23722 14716 23786 14720
rect 23722 14660 23726 14716
rect 23726 14660 23782 14716
rect 23782 14660 23786 14716
rect 23722 14656 23786 14660
rect 23802 14716 23866 14720
rect 23802 14660 23806 14716
rect 23806 14660 23862 14716
rect 23862 14660 23866 14716
rect 23802 14656 23866 14660
rect 23882 14716 23946 14720
rect 23882 14660 23886 14716
rect 23886 14660 23942 14716
rect 23942 14660 23946 14716
rect 23882 14656 23946 14660
rect 23962 14716 24026 14720
rect 23962 14660 23966 14716
rect 23966 14660 24022 14716
rect 24022 14660 24026 14716
rect 23962 14656 24026 14660
rect 31496 14716 31560 14720
rect 31496 14660 31500 14716
rect 31500 14660 31556 14716
rect 31556 14660 31560 14716
rect 31496 14656 31560 14660
rect 31576 14716 31640 14720
rect 31576 14660 31580 14716
rect 31580 14660 31636 14716
rect 31636 14660 31640 14716
rect 31576 14656 31640 14660
rect 31656 14716 31720 14720
rect 31656 14660 31660 14716
rect 31660 14660 31716 14716
rect 31716 14660 31720 14716
rect 31656 14656 31720 14660
rect 31736 14716 31800 14720
rect 31736 14660 31740 14716
rect 31740 14660 31796 14716
rect 31796 14660 31800 14716
rect 31736 14656 31800 14660
rect 4287 14172 4351 14176
rect 4287 14116 4291 14172
rect 4291 14116 4347 14172
rect 4347 14116 4351 14172
rect 4287 14112 4351 14116
rect 4367 14172 4431 14176
rect 4367 14116 4371 14172
rect 4371 14116 4427 14172
rect 4427 14116 4431 14172
rect 4367 14112 4431 14116
rect 4447 14172 4511 14176
rect 4447 14116 4451 14172
rect 4451 14116 4507 14172
rect 4507 14116 4511 14172
rect 4447 14112 4511 14116
rect 4527 14172 4591 14176
rect 4527 14116 4531 14172
rect 4531 14116 4587 14172
rect 4587 14116 4591 14172
rect 4527 14112 4591 14116
rect 12061 14172 12125 14176
rect 12061 14116 12065 14172
rect 12065 14116 12121 14172
rect 12121 14116 12125 14172
rect 12061 14112 12125 14116
rect 12141 14172 12205 14176
rect 12141 14116 12145 14172
rect 12145 14116 12201 14172
rect 12201 14116 12205 14172
rect 12141 14112 12205 14116
rect 12221 14172 12285 14176
rect 12221 14116 12225 14172
rect 12225 14116 12281 14172
rect 12281 14116 12285 14172
rect 12221 14112 12285 14116
rect 12301 14172 12365 14176
rect 12301 14116 12305 14172
rect 12305 14116 12361 14172
rect 12361 14116 12365 14172
rect 12301 14112 12365 14116
rect 19835 14172 19899 14176
rect 19835 14116 19839 14172
rect 19839 14116 19895 14172
rect 19895 14116 19899 14172
rect 19835 14112 19899 14116
rect 19915 14172 19979 14176
rect 19915 14116 19919 14172
rect 19919 14116 19975 14172
rect 19975 14116 19979 14172
rect 19915 14112 19979 14116
rect 19995 14172 20059 14176
rect 19995 14116 19999 14172
rect 19999 14116 20055 14172
rect 20055 14116 20059 14172
rect 19995 14112 20059 14116
rect 20075 14172 20139 14176
rect 20075 14116 20079 14172
rect 20079 14116 20135 14172
rect 20135 14116 20139 14172
rect 20075 14112 20139 14116
rect 27609 14172 27673 14176
rect 27609 14116 27613 14172
rect 27613 14116 27669 14172
rect 27669 14116 27673 14172
rect 27609 14112 27673 14116
rect 27689 14172 27753 14176
rect 27689 14116 27693 14172
rect 27693 14116 27749 14172
rect 27749 14116 27753 14172
rect 27689 14112 27753 14116
rect 27769 14172 27833 14176
rect 27769 14116 27773 14172
rect 27773 14116 27829 14172
rect 27829 14116 27833 14172
rect 27769 14112 27833 14116
rect 27849 14172 27913 14176
rect 27849 14116 27853 14172
rect 27853 14116 27909 14172
rect 27909 14116 27913 14172
rect 27849 14112 27913 14116
rect 8174 13628 8238 13632
rect 8174 13572 8178 13628
rect 8178 13572 8234 13628
rect 8234 13572 8238 13628
rect 8174 13568 8238 13572
rect 8254 13628 8318 13632
rect 8254 13572 8258 13628
rect 8258 13572 8314 13628
rect 8314 13572 8318 13628
rect 8254 13568 8318 13572
rect 8334 13628 8398 13632
rect 8334 13572 8338 13628
rect 8338 13572 8394 13628
rect 8394 13572 8398 13628
rect 8334 13568 8398 13572
rect 8414 13628 8478 13632
rect 8414 13572 8418 13628
rect 8418 13572 8474 13628
rect 8474 13572 8478 13628
rect 8414 13568 8478 13572
rect 15948 13628 16012 13632
rect 15948 13572 15952 13628
rect 15952 13572 16008 13628
rect 16008 13572 16012 13628
rect 15948 13568 16012 13572
rect 16028 13628 16092 13632
rect 16028 13572 16032 13628
rect 16032 13572 16088 13628
rect 16088 13572 16092 13628
rect 16028 13568 16092 13572
rect 16108 13628 16172 13632
rect 16108 13572 16112 13628
rect 16112 13572 16168 13628
rect 16168 13572 16172 13628
rect 16108 13568 16172 13572
rect 16188 13628 16252 13632
rect 16188 13572 16192 13628
rect 16192 13572 16248 13628
rect 16248 13572 16252 13628
rect 16188 13568 16252 13572
rect 23722 13628 23786 13632
rect 23722 13572 23726 13628
rect 23726 13572 23782 13628
rect 23782 13572 23786 13628
rect 23722 13568 23786 13572
rect 23802 13628 23866 13632
rect 23802 13572 23806 13628
rect 23806 13572 23862 13628
rect 23862 13572 23866 13628
rect 23802 13568 23866 13572
rect 23882 13628 23946 13632
rect 23882 13572 23886 13628
rect 23886 13572 23942 13628
rect 23942 13572 23946 13628
rect 23882 13568 23946 13572
rect 23962 13628 24026 13632
rect 23962 13572 23966 13628
rect 23966 13572 24022 13628
rect 24022 13572 24026 13628
rect 23962 13568 24026 13572
rect 31496 13628 31560 13632
rect 31496 13572 31500 13628
rect 31500 13572 31556 13628
rect 31556 13572 31560 13628
rect 31496 13568 31560 13572
rect 31576 13628 31640 13632
rect 31576 13572 31580 13628
rect 31580 13572 31636 13628
rect 31636 13572 31640 13628
rect 31576 13568 31640 13572
rect 31656 13628 31720 13632
rect 31656 13572 31660 13628
rect 31660 13572 31716 13628
rect 31716 13572 31720 13628
rect 31656 13568 31720 13572
rect 31736 13628 31800 13632
rect 31736 13572 31740 13628
rect 31740 13572 31796 13628
rect 31796 13572 31800 13628
rect 31736 13568 31800 13572
rect 4287 13084 4351 13088
rect 4287 13028 4291 13084
rect 4291 13028 4347 13084
rect 4347 13028 4351 13084
rect 4287 13024 4351 13028
rect 4367 13084 4431 13088
rect 4367 13028 4371 13084
rect 4371 13028 4427 13084
rect 4427 13028 4431 13084
rect 4367 13024 4431 13028
rect 4447 13084 4511 13088
rect 4447 13028 4451 13084
rect 4451 13028 4507 13084
rect 4507 13028 4511 13084
rect 4447 13024 4511 13028
rect 4527 13084 4591 13088
rect 4527 13028 4531 13084
rect 4531 13028 4587 13084
rect 4587 13028 4591 13084
rect 4527 13024 4591 13028
rect 12061 13084 12125 13088
rect 12061 13028 12065 13084
rect 12065 13028 12121 13084
rect 12121 13028 12125 13084
rect 12061 13024 12125 13028
rect 12141 13084 12205 13088
rect 12141 13028 12145 13084
rect 12145 13028 12201 13084
rect 12201 13028 12205 13084
rect 12141 13024 12205 13028
rect 12221 13084 12285 13088
rect 12221 13028 12225 13084
rect 12225 13028 12281 13084
rect 12281 13028 12285 13084
rect 12221 13024 12285 13028
rect 12301 13084 12365 13088
rect 12301 13028 12305 13084
rect 12305 13028 12361 13084
rect 12361 13028 12365 13084
rect 12301 13024 12365 13028
rect 19835 13084 19899 13088
rect 19835 13028 19839 13084
rect 19839 13028 19895 13084
rect 19895 13028 19899 13084
rect 19835 13024 19899 13028
rect 19915 13084 19979 13088
rect 19915 13028 19919 13084
rect 19919 13028 19975 13084
rect 19975 13028 19979 13084
rect 19915 13024 19979 13028
rect 19995 13084 20059 13088
rect 19995 13028 19999 13084
rect 19999 13028 20055 13084
rect 20055 13028 20059 13084
rect 19995 13024 20059 13028
rect 20075 13084 20139 13088
rect 20075 13028 20079 13084
rect 20079 13028 20135 13084
rect 20135 13028 20139 13084
rect 20075 13024 20139 13028
rect 27609 13084 27673 13088
rect 27609 13028 27613 13084
rect 27613 13028 27669 13084
rect 27669 13028 27673 13084
rect 27609 13024 27673 13028
rect 27689 13084 27753 13088
rect 27689 13028 27693 13084
rect 27693 13028 27749 13084
rect 27749 13028 27753 13084
rect 27689 13024 27753 13028
rect 27769 13084 27833 13088
rect 27769 13028 27773 13084
rect 27773 13028 27829 13084
rect 27829 13028 27833 13084
rect 27769 13024 27833 13028
rect 27849 13084 27913 13088
rect 27849 13028 27853 13084
rect 27853 13028 27909 13084
rect 27909 13028 27913 13084
rect 27849 13024 27913 13028
rect 8174 12540 8238 12544
rect 8174 12484 8178 12540
rect 8178 12484 8234 12540
rect 8234 12484 8238 12540
rect 8174 12480 8238 12484
rect 8254 12540 8318 12544
rect 8254 12484 8258 12540
rect 8258 12484 8314 12540
rect 8314 12484 8318 12540
rect 8254 12480 8318 12484
rect 8334 12540 8398 12544
rect 8334 12484 8338 12540
rect 8338 12484 8394 12540
rect 8394 12484 8398 12540
rect 8334 12480 8398 12484
rect 8414 12540 8478 12544
rect 8414 12484 8418 12540
rect 8418 12484 8474 12540
rect 8474 12484 8478 12540
rect 8414 12480 8478 12484
rect 15948 12540 16012 12544
rect 15948 12484 15952 12540
rect 15952 12484 16008 12540
rect 16008 12484 16012 12540
rect 15948 12480 16012 12484
rect 16028 12540 16092 12544
rect 16028 12484 16032 12540
rect 16032 12484 16088 12540
rect 16088 12484 16092 12540
rect 16028 12480 16092 12484
rect 16108 12540 16172 12544
rect 16108 12484 16112 12540
rect 16112 12484 16168 12540
rect 16168 12484 16172 12540
rect 16108 12480 16172 12484
rect 16188 12540 16252 12544
rect 16188 12484 16192 12540
rect 16192 12484 16248 12540
rect 16248 12484 16252 12540
rect 16188 12480 16252 12484
rect 23722 12540 23786 12544
rect 23722 12484 23726 12540
rect 23726 12484 23782 12540
rect 23782 12484 23786 12540
rect 23722 12480 23786 12484
rect 23802 12540 23866 12544
rect 23802 12484 23806 12540
rect 23806 12484 23862 12540
rect 23862 12484 23866 12540
rect 23802 12480 23866 12484
rect 23882 12540 23946 12544
rect 23882 12484 23886 12540
rect 23886 12484 23942 12540
rect 23942 12484 23946 12540
rect 23882 12480 23946 12484
rect 23962 12540 24026 12544
rect 23962 12484 23966 12540
rect 23966 12484 24022 12540
rect 24022 12484 24026 12540
rect 23962 12480 24026 12484
rect 31496 12540 31560 12544
rect 31496 12484 31500 12540
rect 31500 12484 31556 12540
rect 31556 12484 31560 12540
rect 31496 12480 31560 12484
rect 31576 12540 31640 12544
rect 31576 12484 31580 12540
rect 31580 12484 31636 12540
rect 31636 12484 31640 12540
rect 31576 12480 31640 12484
rect 31656 12540 31720 12544
rect 31656 12484 31660 12540
rect 31660 12484 31716 12540
rect 31716 12484 31720 12540
rect 31656 12480 31720 12484
rect 31736 12540 31800 12544
rect 31736 12484 31740 12540
rect 31740 12484 31796 12540
rect 31796 12484 31800 12540
rect 31736 12480 31800 12484
rect 4287 11996 4351 12000
rect 4287 11940 4291 11996
rect 4291 11940 4347 11996
rect 4347 11940 4351 11996
rect 4287 11936 4351 11940
rect 4367 11996 4431 12000
rect 4367 11940 4371 11996
rect 4371 11940 4427 11996
rect 4427 11940 4431 11996
rect 4367 11936 4431 11940
rect 4447 11996 4511 12000
rect 4447 11940 4451 11996
rect 4451 11940 4507 11996
rect 4507 11940 4511 11996
rect 4447 11936 4511 11940
rect 4527 11996 4591 12000
rect 4527 11940 4531 11996
rect 4531 11940 4587 11996
rect 4587 11940 4591 11996
rect 4527 11936 4591 11940
rect 12061 11996 12125 12000
rect 12061 11940 12065 11996
rect 12065 11940 12121 11996
rect 12121 11940 12125 11996
rect 12061 11936 12125 11940
rect 12141 11996 12205 12000
rect 12141 11940 12145 11996
rect 12145 11940 12201 11996
rect 12201 11940 12205 11996
rect 12141 11936 12205 11940
rect 12221 11996 12285 12000
rect 12221 11940 12225 11996
rect 12225 11940 12281 11996
rect 12281 11940 12285 11996
rect 12221 11936 12285 11940
rect 12301 11996 12365 12000
rect 12301 11940 12305 11996
rect 12305 11940 12361 11996
rect 12361 11940 12365 11996
rect 12301 11936 12365 11940
rect 19835 11996 19899 12000
rect 19835 11940 19839 11996
rect 19839 11940 19895 11996
rect 19895 11940 19899 11996
rect 19835 11936 19899 11940
rect 19915 11996 19979 12000
rect 19915 11940 19919 11996
rect 19919 11940 19975 11996
rect 19975 11940 19979 11996
rect 19915 11936 19979 11940
rect 19995 11996 20059 12000
rect 19995 11940 19999 11996
rect 19999 11940 20055 11996
rect 20055 11940 20059 11996
rect 19995 11936 20059 11940
rect 20075 11996 20139 12000
rect 20075 11940 20079 11996
rect 20079 11940 20135 11996
rect 20135 11940 20139 11996
rect 20075 11936 20139 11940
rect 27609 11996 27673 12000
rect 27609 11940 27613 11996
rect 27613 11940 27669 11996
rect 27669 11940 27673 11996
rect 27609 11936 27673 11940
rect 27689 11996 27753 12000
rect 27689 11940 27693 11996
rect 27693 11940 27749 11996
rect 27749 11940 27753 11996
rect 27689 11936 27753 11940
rect 27769 11996 27833 12000
rect 27769 11940 27773 11996
rect 27773 11940 27829 11996
rect 27829 11940 27833 11996
rect 27769 11936 27833 11940
rect 27849 11996 27913 12000
rect 27849 11940 27853 11996
rect 27853 11940 27909 11996
rect 27909 11940 27913 11996
rect 27849 11936 27913 11940
rect 8174 11452 8238 11456
rect 8174 11396 8178 11452
rect 8178 11396 8234 11452
rect 8234 11396 8238 11452
rect 8174 11392 8238 11396
rect 8254 11452 8318 11456
rect 8254 11396 8258 11452
rect 8258 11396 8314 11452
rect 8314 11396 8318 11452
rect 8254 11392 8318 11396
rect 8334 11452 8398 11456
rect 8334 11396 8338 11452
rect 8338 11396 8394 11452
rect 8394 11396 8398 11452
rect 8334 11392 8398 11396
rect 8414 11452 8478 11456
rect 8414 11396 8418 11452
rect 8418 11396 8474 11452
rect 8474 11396 8478 11452
rect 8414 11392 8478 11396
rect 15948 11452 16012 11456
rect 15948 11396 15952 11452
rect 15952 11396 16008 11452
rect 16008 11396 16012 11452
rect 15948 11392 16012 11396
rect 16028 11452 16092 11456
rect 16028 11396 16032 11452
rect 16032 11396 16088 11452
rect 16088 11396 16092 11452
rect 16028 11392 16092 11396
rect 16108 11452 16172 11456
rect 16108 11396 16112 11452
rect 16112 11396 16168 11452
rect 16168 11396 16172 11452
rect 16108 11392 16172 11396
rect 16188 11452 16252 11456
rect 16188 11396 16192 11452
rect 16192 11396 16248 11452
rect 16248 11396 16252 11452
rect 16188 11392 16252 11396
rect 23722 11452 23786 11456
rect 23722 11396 23726 11452
rect 23726 11396 23782 11452
rect 23782 11396 23786 11452
rect 23722 11392 23786 11396
rect 23802 11452 23866 11456
rect 23802 11396 23806 11452
rect 23806 11396 23862 11452
rect 23862 11396 23866 11452
rect 23802 11392 23866 11396
rect 23882 11452 23946 11456
rect 23882 11396 23886 11452
rect 23886 11396 23942 11452
rect 23942 11396 23946 11452
rect 23882 11392 23946 11396
rect 23962 11452 24026 11456
rect 23962 11396 23966 11452
rect 23966 11396 24022 11452
rect 24022 11396 24026 11452
rect 23962 11392 24026 11396
rect 31496 11452 31560 11456
rect 31496 11396 31500 11452
rect 31500 11396 31556 11452
rect 31556 11396 31560 11452
rect 31496 11392 31560 11396
rect 31576 11452 31640 11456
rect 31576 11396 31580 11452
rect 31580 11396 31636 11452
rect 31636 11396 31640 11452
rect 31576 11392 31640 11396
rect 31656 11452 31720 11456
rect 31656 11396 31660 11452
rect 31660 11396 31716 11452
rect 31716 11396 31720 11452
rect 31656 11392 31720 11396
rect 31736 11452 31800 11456
rect 31736 11396 31740 11452
rect 31740 11396 31796 11452
rect 31796 11396 31800 11452
rect 31736 11392 31800 11396
rect 4287 10908 4351 10912
rect 4287 10852 4291 10908
rect 4291 10852 4347 10908
rect 4347 10852 4351 10908
rect 4287 10848 4351 10852
rect 4367 10908 4431 10912
rect 4367 10852 4371 10908
rect 4371 10852 4427 10908
rect 4427 10852 4431 10908
rect 4367 10848 4431 10852
rect 4447 10908 4511 10912
rect 4447 10852 4451 10908
rect 4451 10852 4507 10908
rect 4507 10852 4511 10908
rect 4447 10848 4511 10852
rect 4527 10908 4591 10912
rect 4527 10852 4531 10908
rect 4531 10852 4587 10908
rect 4587 10852 4591 10908
rect 4527 10848 4591 10852
rect 12061 10908 12125 10912
rect 12061 10852 12065 10908
rect 12065 10852 12121 10908
rect 12121 10852 12125 10908
rect 12061 10848 12125 10852
rect 12141 10908 12205 10912
rect 12141 10852 12145 10908
rect 12145 10852 12201 10908
rect 12201 10852 12205 10908
rect 12141 10848 12205 10852
rect 12221 10908 12285 10912
rect 12221 10852 12225 10908
rect 12225 10852 12281 10908
rect 12281 10852 12285 10908
rect 12221 10848 12285 10852
rect 12301 10908 12365 10912
rect 12301 10852 12305 10908
rect 12305 10852 12361 10908
rect 12361 10852 12365 10908
rect 12301 10848 12365 10852
rect 19835 10908 19899 10912
rect 19835 10852 19839 10908
rect 19839 10852 19895 10908
rect 19895 10852 19899 10908
rect 19835 10848 19899 10852
rect 19915 10908 19979 10912
rect 19915 10852 19919 10908
rect 19919 10852 19975 10908
rect 19975 10852 19979 10908
rect 19915 10848 19979 10852
rect 19995 10908 20059 10912
rect 19995 10852 19999 10908
rect 19999 10852 20055 10908
rect 20055 10852 20059 10908
rect 19995 10848 20059 10852
rect 20075 10908 20139 10912
rect 20075 10852 20079 10908
rect 20079 10852 20135 10908
rect 20135 10852 20139 10908
rect 20075 10848 20139 10852
rect 27609 10908 27673 10912
rect 27609 10852 27613 10908
rect 27613 10852 27669 10908
rect 27669 10852 27673 10908
rect 27609 10848 27673 10852
rect 27689 10908 27753 10912
rect 27689 10852 27693 10908
rect 27693 10852 27749 10908
rect 27749 10852 27753 10908
rect 27689 10848 27753 10852
rect 27769 10908 27833 10912
rect 27769 10852 27773 10908
rect 27773 10852 27829 10908
rect 27829 10852 27833 10908
rect 27769 10848 27833 10852
rect 27849 10908 27913 10912
rect 27849 10852 27853 10908
rect 27853 10852 27909 10908
rect 27909 10852 27913 10908
rect 27849 10848 27913 10852
rect 8174 10364 8238 10368
rect 8174 10308 8178 10364
rect 8178 10308 8234 10364
rect 8234 10308 8238 10364
rect 8174 10304 8238 10308
rect 8254 10364 8318 10368
rect 8254 10308 8258 10364
rect 8258 10308 8314 10364
rect 8314 10308 8318 10364
rect 8254 10304 8318 10308
rect 8334 10364 8398 10368
rect 8334 10308 8338 10364
rect 8338 10308 8394 10364
rect 8394 10308 8398 10364
rect 8334 10304 8398 10308
rect 8414 10364 8478 10368
rect 8414 10308 8418 10364
rect 8418 10308 8474 10364
rect 8474 10308 8478 10364
rect 8414 10304 8478 10308
rect 15948 10364 16012 10368
rect 15948 10308 15952 10364
rect 15952 10308 16008 10364
rect 16008 10308 16012 10364
rect 15948 10304 16012 10308
rect 16028 10364 16092 10368
rect 16028 10308 16032 10364
rect 16032 10308 16088 10364
rect 16088 10308 16092 10364
rect 16028 10304 16092 10308
rect 16108 10364 16172 10368
rect 16108 10308 16112 10364
rect 16112 10308 16168 10364
rect 16168 10308 16172 10364
rect 16108 10304 16172 10308
rect 16188 10364 16252 10368
rect 16188 10308 16192 10364
rect 16192 10308 16248 10364
rect 16248 10308 16252 10364
rect 16188 10304 16252 10308
rect 23722 10364 23786 10368
rect 23722 10308 23726 10364
rect 23726 10308 23782 10364
rect 23782 10308 23786 10364
rect 23722 10304 23786 10308
rect 23802 10364 23866 10368
rect 23802 10308 23806 10364
rect 23806 10308 23862 10364
rect 23862 10308 23866 10364
rect 23802 10304 23866 10308
rect 23882 10364 23946 10368
rect 23882 10308 23886 10364
rect 23886 10308 23942 10364
rect 23942 10308 23946 10364
rect 23882 10304 23946 10308
rect 23962 10364 24026 10368
rect 23962 10308 23966 10364
rect 23966 10308 24022 10364
rect 24022 10308 24026 10364
rect 23962 10304 24026 10308
rect 31496 10364 31560 10368
rect 31496 10308 31500 10364
rect 31500 10308 31556 10364
rect 31556 10308 31560 10364
rect 31496 10304 31560 10308
rect 31576 10364 31640 10368
rect 31576 10308 31580 10364
rect 31580 10308 31636 10364
rect 31636 10308 31640 10364
rect 31576 10304 31640 10308
rect 31656 10364 31720 10368
rect 31656 10308 31660 10364
rect 31660 10308 31716 10364
rect 31716 10308 31720 10364
rect 31656 10304 31720 10308
rect 31736 10364 31800 10368
rect 31736 10308 31740 10364
rect 31740 10308 31796 10364
rect 31796 10308 31800 10364
rect 31736 10304 31800 10308
rect 4287 9820 4351 9824
rect 4287 9764 4291 9820
rect 4291 9764 4347 9820
rect 4347 9764 4351 9820
rect 4287 9760 4351 9764
rect 4367 9820 4431 9824
rect 4367 9764 4371 9820
rect 4371 9764 4427 9820
rect 4427 9764 4431 9820
rect 4367 9760 4431 9764
rect 4447 9820 4511 9824
rect 4447 9764 4451 9820
rect 4451 9764 4507 9820
rect 4507 9764 4511 9820
rect 4447 9760 4511 9764
rect 4527 9820 4591 9824
rect 4527 9764 4531 9820
rect 4531 9764 4587 9820
rect 4587 9764 4591 9820
rect 4527 9760 4591 9764
rect 12061 9820 12125 9824
rect 12061 9764 12065 9820
rect 12065 9764 12121 9820
rect 12121 9764 12125 9820
rect 12061 9760 12125 9764
rect 12141 9820 12205 9824
rect 12141 9764 12145 9820
rect 12145 9764 12201 9820
rect 12201 9764 12205 9820
rect 12141 9760 12205 9764
rect 12221 9820 12285 9824
rect 12221 9764 12225 9820
rect 12225 9764 12281 9820
rect 12281 9764 12285 9820
rect 12221 9760 12285 9764
rect 12301 9820 12365 9824
rect 12301 9764 12305 9820
rect 12305 9764 12361 9820
rect 12361 9764 12365 9820
rect 12301 9760 12365 9764
rect 19835 9820 19899 9824
rect 19835 9764 19839 9820
rect 19839 9764 19895 9820
rect 19895 9764 19899 9820
rect 19835 9760 19899 9764
rect 19915 9820 19979 9824
rect 19915 9764 19919 9820
rect 19919 9764 19975 9820
rect 19975 9764 19979 9820
rect 19915 9760 19979 9764
rect 19995 9820 20059 9824
rect 19995 9764 19999 9820
rect 19999 9764 20055 9820
rect 20055 9764 20059 9820
rect 19995 9760 20059 9764
rect 20075 9820 20139 9824
rect 20075 9764 20079 9820
rect 20079 9764 20135 9820
rect 20135 9764 20139 9820
rect 20075 9760 20139 9764
rect 27609 9820 27673 9824
rect 27609 9764 27613 9820
rect 27613 9764 27669 9820
rect 27669 9764 27673 9820
rect 27609 9760 27673 9764
rect 27689 9820 27753 9824
rect 27689 9764 27693 9820
rect 27693 9764 27749 9820
rect 27749 9764 27753 9820
rect 27689 9760 27753 9764
rect 27769 9820 27833 9824
rect 27769 9764 27773 9820
rect 27773 9764 27829 9820
rect 27829 9764 27833 9820
rect 27769 9760 27833 9764
rect 27849 9820 27913 9824
rect 27849 9764 27853 9820
rect 27853 9764 27909 9820
rect 27909 9764 27913 9820
rect 27849 9760 27913 9764
rect 8174 9276 8238 9280
rect 8174 9220 8178 9276
rect 8178 9220 8234 9276
rect 8234 9220 8238 9276
rect 8174 9216 8238 9220
rect 8254 9276 8318 9280
rect 8254 9220 8258 9276
rect 8258 9220 8314 9276
rect 8314 9220 8318 9276
rect 8254 9216 8318 9220
rect 8334 9276 8398 9280
rect 8334 9220 8338 9276
rect 8338 9220 8394 9276
rect 8394 9220 8398 9276
rect 8334 9216 8398 9220
rect 8414 9276 8478 9280
rect 8414 9220 8418 9276
rect 8418 9220 8474 9276
rect 8474 9220 8478 9276
rect 8414 9216 8478 9220
rect 15948 9276 16012 9280
rect 15948 9220 15952 9276
rect 15952 9220 16008 9276
rect 16008 9220 16012 9276
rect 15948 9216 16012 9220
rect 16028 9276 16092 9280
rect 16028 9220 16032 9276
rect 16032 9220 16088 9276
rect 16088 9220 16092 9276
rect 16028 9216 16092 9220
rect 16108 9276 16172 9280
rect 16108 9220 16112 9276
rect 16112 9220 16168 9276
rect 16168 9220 16172 9276
rect 16108 9216 16172 9220
rect 16188 9276 16252 9280
rect 16188 9220 16192 9276
rect 16192 9220 16248 9276
rect 16248 9220 16252 9276
rect 16188 9216 16252 9220
rect 23722 9276 23786 9280
rect 23722 9220 23726 9276
rect 23726 9220 23782 9276
rect 23782 9220 23786 9276
rect 23722 9216 23786 9220
rect 23802 9276 23866 9280
rect 23802 9220 23806 9276
rect 23806 9220 23862 9276
rect 23862 9220 23866 9276
rect 23802 9216 23866 9220
rect 23882 9276 23946 9280
rect 23882 9220 23886 9276
rect 23886 9220 23942 9276
rect 23942 9220 23946 9276
rect 23882 9216 23946 9220
rect 23962 9276 24026 9280
rect 23962 9220 23966 9276
rect 23966 9220 24022 9276
rect 24022 9220 24026 9276
rect 23962 9216 24026 9220
rect 31496 9276 31560 9280
rect 31496 9220 31500 9276
rect 31500 9220 31556 9276
rect 31556 9220 31560 9276
rect 31496 9216 31560 9220
rect 31576 9276 31640 9280
rect 31576 9220 31580 9276
rect 31580 9220 31636 9276
rect 31636 9220 31640 9276
rect 31576 9216 31640 9220
rect 31656 9276 31720 9280
rect 31656 9220 31660 9276
rect 31660 9220 31716 9276
rect 31716 9220 31720 9276
rect 31656 9216 31720 9220
rect 31736 9276 31800 9280
rect 31736 9220 31740 9276
rect 31740 9220 31796 9276
rect 31796 9220 31800 9276
rect 31736 9216 31800 9220
rect 4287 8732 4351 8736
rect 4287 8676 4291 8732
rect 4291 8676 4347 8732
rect 4347 8676 4351 8732
rect 4287 8672 4351 8676
rect 4367 8732 4431 8736
rect 4367 8676 4371 8732
rect 4371 8676 4427 8732
rect 4427 8676 4431 8732
rect 4367 8672 4431 8676
rect 4447 8732 4511 8736
rect 4447 8676 4451 8732
rect 4451 8676 4507 8732
rect 4507 8676 4511 8732
rect 4447 8672 4511 8676
rect 4527 8732 4591 8736
rect 4527 8676 4531 8732
rect 4531 8676 4587 8732
rect 4587 8676 4591 8732
rect 4527 8672 4591 8676
rect 12061 8732 12125 8736
rect 12061 8676 12065 8732
rect 12065 8676 12121 8732
rect 12121 8676 12125 8732
rect 12061 8672 12125 8676
rect 12141 8732 12205 8736
rect 12141 8676 12145 8732
rect 12145 8676 12201 8732
rect 12201 8676 12205 8732
rect 12141 8672 12205 8676
rect 12221 8732 12285 8736
rect 12221 8676 12225 8732
rect 12225 8676 12281 8732
rect 12281 8676 12285 8732
rect 12221 8672 12285 8676
rect 12301 8732 12365 8736
rect 12301 8676 12305 8732
rect 12305 8676 12361 8732
rect 12361 8676 12365 8732
rect 12301 8672 12365 8676
rect 19835 8732 19899 8736
rect 19835 8676 19839 8732
rect 19839 8676 19895 8732
rect 19895 8676 19899 8732
rect 19835 8672 19899 8676
rect 19915 8732 19979 8736
rect 19915 8676 19919 8732
rect 19919 8676 19975 8732
rect 19975 8676 19979 8732
rect 19915 8672 19979 8676
rect 19995 8732 20059 8736
rect 19995 8676 19999 8732
rect 19999 8676 20055 8732
rect 20055 8676 20059 8732
rect 19995 8672 20059 8676
rect 20075 8732 20139 8736
rect 20075 8676 20079 8732
rect 20079 8676 20135 8732
rect 20135 8676 20139 8732
rect 20075 8672 20139 8676
rect 27609 8732 27673 8736
rect 27609 8676 27613 8732
rect 27613 8676 27669 8732
rect 27669 8676 27673 8732
rect 27609 8672 27673 8676
rect 27689 8732 27753 8736
rect 27689 8676 27693 8732
rect 27693 8676 27749 8732
rect 27749 8676 27753 8732
rect 27689 8672 27753 8676
rect 27769 8732 27833 8736
rect 27769 8676 27773 8732
rect 27773 8676 27829 8732
rect 27829 8676 27833 8732
rect 27769 8672 27833 8676
rect 27849 8732 27913 8736
rect 27849 8676 27853 8732
rect 27853 8676 27909 8732
rect 27909 8676 27913 8732
rect 27849 8672 27913 8676
rect 8174 8188 8238 8192
rect 8174 8132 8178 8188
rect 8178 8132 8234 8188
rect 8234 8132 8238 8188
rect 8174 8128 8238 8132
rect 8254 8188 8318 8192
rect 8254 8132 8258 8188
rect 8258 8132 8314 8188
rect 8314 8132 8318 8188
rect 8254 8128 8318 8132
rect 8334 8188 8398 8192
rect 8334 8132 8338 8188
rect 8338 8132 8394 8188
rect 8394 8132 8398 8188
rect 8334 8128 8398 8132
rect 8414 8188 8478 8192
rect 8414 8132 8418 8188
rect 8418 8132 8474 8188
rect 8474 8132 8478 8188
rect 8414 8128 8478 8132
rect 15948 8188 16012 8192
rect 15948 8132 15952 8188
rect 15952 8132 16008 8188
rect 16008 8132 16012 8188
rect 15948 8128 16012 8132
rect 16028 8188 16092 8192
rect 16028 8132 16032 8188
rect 16032 8132 16088 8188
rect 16088 8132 16092 8188
rect 16028 8128 16092 8132
rect 16108 8188 16172 8192
rect 16108 8132 16112 8188
rect 16112 8132 16168 8188
rect 16168 8132 16172 8188
rect 16108 8128 16172 8132
rect 16188 8188 16252 8192
rect 16188 8132 16192 8188
rect 16192 8132 16248 8188
rect 16248 8132 16252 8188
rect 16188 8128 16252 8132
rect 23722 8188 23786 8192
rect 23722 8132 23726 8188
rect 23726 8132 23782 8188
rect 23782 8132 23786 8188
rect 23722 8128 23786 8132
rect 23802 8188 23866 8192
rect 23802 8132 23806 8188
rect 23806 8132 23862 8188
rect 23862 8132 23866 8188
rect 23802 8128 23866 8132
rect 23882 8188 23946 8192
rect 23882 8132 23886 8188
rect 23886 8132 23942 8188
rect 23942 8132 23946 8188
rect 23882 8128 23946 8132
rect 23962 8188 24026 8192
rect 23962 8132 23966 8188
rect 23966 8132 24022 8188
rect 24022 8132 24026 8188
rect 23962 8128 24026 8132
rect 31496 8188 31560 8192
rect 31496 8132 31500 8188
rect 31500 8132 31556 8188
rect 31556 8132 31560 8188
rect 31496 8128 31560 8132
rect 31576 8188 31640 8192
rect 31576 8132 31580 8188
rect 31580 8132 31636 8188
rect 31636 8132 31640 8188
rect 31576 8128 31640 8132
rect 31656 8188 31720 8192
rect 31656 8132 31660 8188
rect 31660 8132 31716 8188
rect 31716 8132 31720 8188
rect 31656 8128 31720 8132
rect 31736 8188 31800 8192
rect 31736 8132 31740 8188
rect 31740 8132 31796 8188
rect 31796 8132 31800 8188
rect 31736 8128 31800 8132
rect 4287 7644 4351 7648
rect 4287 7588 4291 7644
rect 4291 7588 4347 7644
rect 4347 7588 4351 7644
rect 4287 7584 4351 7588
rect 4367 7644 4431 7648
rect 4367 7588 4371 7644
rect 4371 7588 4427 7644
rect 4427 7588 4431 7644
rect 4367 7584 4431 7588
rect 4447 7644 4511 7648
rect 4447 7588 4451 7644
rect 4451 7588 4507 7644
rect 4507 7588 4511 7644
rect 4447 7584 4511 7588
rect 4527 7644 4591 7648
rect 4527 7588 4531 7644
rect 4531 7588 4587 7644
rect 4587 7588 4591 7644
rect 4527 7584 4591 7588
rect 12061 7644 12125 7648
rect 12061 7588 12065 7644
rect 12065 7588 12121 7644
rect 12121 7588 12125 7644
rect 12061 7584 12125 7588
rect 12141 7644 12205 7648
rect 12141 7588 12145 7644
rect 12145 7588 12201 7644
rect 12201 7588 12205 7644
rect 12141 7584 12205 7588
rect 12221 7644 12285 7648
rect 12221 7588 12225 7644
rect 12225 7588 12281 7644
rect 12281 7588 12285 7644
rect 12221 7584 12285 7588
rect 12301 7644 12365 7648
rect 12301 7588 12305 7644
rect 12305 7588 12361 7644
rect 12361 7588 12365 7644
rect 12301 7584 12365 7588
rect 19835 7644 19899 7648
rect 19835 7588 19839 7644
rect 19839 7588 19895 7644
rect 19895 7588 19899 7644
rect 19835 7584 19899 7588
rect 19915 7644 19979 7648
rect 19915 7588 19919 7644
rect 19919 7588 19975 7644
rect 19975 7588 19979 7644
rect 19915 7584 19979 7588
rect 19995 7644 20059 7648
rect 19995 7588 19999 7644
rect 19999 7588 20055 7644
rect 20055 7588 20059 7644
rect 19995 7584 20059 7588
rect 20075 7644 20139 7648
rect 20075 7588 20079 7644
rect 20079 7588 20135 7644
rect 20135 7588 20139 7644
rect 20075 7584 20139 7588
rect 27609 7644 27673 7648
rect 27609 7588 27613 7644
rect 27613 7588 27669 7644
rect 27669 7588 27673 7644
rect 27609 7584 27673 7588
rect 27689 7644 27753 7648
rect 27689 7588 27693 7644
rect 27693 7588 27749 7644
rect 27749 7588 27753 7644
rect 27689 7584 27753 7588
rect 27769 7644 27833 7648
rect 27769 7588 27773 7644
rect 27773 7588 27829 7644
rect 27829 7588 27833 7644
rect 27769 7584 27833 7588
rect 27849 7644 27913 7648
rect 27849 7588 27853 7644
rect 27853 7588 27909 7644
rect 27909 7588 27913 7644
rect 27849 7584 27913 7588
rect 8174 7100 8238 7104
rect 8174 7044 8178 7100
rect 8178 7044 8234 7100
rect 8234 7044 8238 7100
rect 8174 7040 8238 7044
rect 8254 7100 8318 7104
rect 8254 7044 8258 7100
rect 8258 7044 8314 7100
rect 8314 7044 8318 7100
rect 8254 7040 8318 7044
rect 8334 7100 8398 7104
rect 8334 7044 8338 7100
rect 8338 7044 8394 7100
rect 8394 7044 8398 7100
rect 8334 7040 8398 7044
rect 8414 7100 8478 7104
rect 8414 7044 8418 7100
rect 8418 7044 8474 7100
rect 8474 7044 8478 7100
rect 8414 7040 8478 7044
rect 15948 7100 16012 7104
rect 15948 7044 15952 7100
rect 15952 7044 16008 7100
rect 16008 7044 16012 7100
rect 15948 7040 16012 7044
rect 16028 7100 16092 7104
rect 16028 7044 16032 7100
rect 16032 7044 16088 7100
rect 16088 7044 16092 7100
rect 16028 7040 16092 7044
rect 16108 7100 16172 7104
rect 16108 7044 16112 7100
rect 16112 7044 16168 7100
rect 16168 7044 16172 7100
rect 16108 7040 16172 7044
rect 16188 7100 16252 7104
rect 16188 7044 16192 7100
rect 16192 7044 16248 7100
rect 16248 7044 16252 7100
rect 16188 7040 16252 7044
rect 23722 7100 23786 7104
rect 23722 7044 23726 7100
rect 23726 7044 23782 7100
rect 23782 7044 23786 7100
rect 23722 7040 23786 7044
rect 23802 7100 23866 7104
rect 23802 7044 23806 7100
rect 23806 7044 23862 7100
rect 23862 7044 23866 7100
rect 23802 7040 23866 7044
rect 23882 7100 23946 7104
rect 23882 7044 23886 7100
rect 23886 7044 23942 7100
rect 23942 7044 23946 7100
rect 23882 7040 23946 7044
rect 23962 7100 24026 7104
rect 23962 7044 23966 7100
rect 23966 7044 24022 7100
rect 24022 7044 24026 7100
rect 23962 7040 24026 7044
rect 31496 7100 31560 7104
rect 31496 7044 31500 7100
rect 31500 7044 31556 7100
rect 31556 7044 31560 7100
rect 31496 7040 31560 7044
rect 31576 7100 31640 7104
rect 31576 7044 31580 7100
rect 31580 7044 31636 7100
rect 31636 7044 31640 7100
rect 31576 7040 31640 7044
rect 31656 7100 31720 7104
rect 31656 7044 31660 7100
rect 31660 7044 31716 7100
rect 31716 7044 31720 7100
rect 31656 7040 31720 7044
rect 31736 7100 31800 7104
rect 31736 7044 31740 7100
rect 31740 7044 31796 7100
rect 31796 7044 31800 7100
rect 31736 7040 31800 7044
rect 4287 6556 4351 6560
rect 4287 6500 4291 6556
rect 4291 6500 4347 6556
rect 4347 6500 4351 6556
rect 4287 6496 4351 6500
rect 4367 6556 4431 6560
rect 4367 6500 4371 6556
rect 4371 6500 4427 6556
rect 4427 6500 4431 6556
rect 4367 6496 4431 6500
rect 4447 6556 4511 6560
rect 4447 6500 4451 6556
rect 4451 6500 4507 6556
rect 4507 6500 4511 6556
rect 4447 6496 4511 6500
rect 4527 6556 4591 6560
rect 4527 6500 4531 6556
rect 4531 6500 4587 6556
rect 4587 6500 4591 6556
rect 4527 6496 4591 6500
rect 12061 6556 12125 6560
rect 12061 6500 12065 6556
rect 12065 6500 12121 6556
rect 12121 6500 12125 6556
rect 12061 6496 12125 6500
rect 12141 6556 12205 6560
rect 12141 6500 12145 6556
rect 12145 6500 12201 6556
rect 12201 6500 12205 6556
rect 12141 6496 12205 6500
rect 12221 6556 12285 6560
rect 12221 6500 12225 6556
rect 12225 6500 12281 6556
rect 12281 6500 12285 6556
rect 12221 6496 12285 6500
rect 12301 6556 12365 6560
rect 12301 6500 12305 6556
rect 12305 6500 12361 6556
rect 12361 6500 12365 6556
rect 12301 6496 12365 6500
rect 19835 6556 19899 6560
rect 19835 6500 19839 6556
rect 19839 6500 19895 6556
rect 19895 6500 19899 6556
rect 19835 6496 19899 6500
rect 19915 6556 19979 6560
rect 19915 6500 19919 6556
rect 19919 6500 19975 6556
rect 19975 6500 19979 6556
rect 19915 6496 19979 6500
rect 19995 6556 20059 6560
rect 19995 6500 19999 6556
rect 19999 6500 20055 6556
rect 20055 6500 20059 6556
rect 19995 6496 20059 6500
rect 20075 6556 20139 6560
rect 20075 6500 20079 6556
rect 20079 6500 20135 6556
rect 20135 6500 20139 6556
rect 20075 6496 20139 6500
rect 27609 6556 27673 6560
rect 27609 6500 27613 6556
rect 27613 6500 27669 6556
rect 27669 6500 27673 6556
rect 27609 6496 27673 6500
rect 27689 6556 27753 6560
rect 27689 6500 27693 6556
rect 27693 6500 27749 6556
rect 27749 6500 27753 6556
rect 27689 6496 27753 6500
rect 27769 6556 27833 6560
rect 27769 6500 27773 6556
rect 27773 6500 27829 6556
rect 27829 6500 27833 6556
rect 27769 6496 27833 6500
rect 27849 6556 27913 6560
rect 27849 6500 27853 6556
rect 27853 6500 27909 6556
rect 27909 6500 27913 6556
rect 27849 6496 27913 6500
rect 8174 6012 8238 6016
rect 8174 5956 8178 6012
rect 8178 5956 8234 6012
rect 8234 5956 8238 6012
rect 8174 5952 8238 5956
rect 8254 6012 8318 6016
rect 8254 5956 8258 6012
rect 8258 5956 8314 6012
rect 8314 5956 8318 6012
rect 8254 5952 8318 5956
rect 8334 6012 8398 6016
rect 8334 5956 8338 6012
rect 8338 5956 8394 6012
rect 8394 5956 8398 6012
rect 8334 5952 8398 5956
rect 8414 6012 8478 6016
rect 8414 5956 8418 6012
rect 8418 5956 8474 6012
rect 8474 5956 8478 6012
rect 8414 5952 8478 5956
rect 15948 6012 16012 6016
rect 15948 5956 15952 6012
rect 15952 5956 16008 6012
rect 16008 5956 16012 6012
rect 15948 5952 16012 5956
rect 16028 6012 16092 6016
rect 16028 5956 16032 6012
rect 16032 5956 16088 6012
rect 16088 5956 16092 6012
rect 16028 5952 16092 5956
rect 16108 6012 16172 6016
rect 16108 5956 16112 6012
rect 16112 5956 16168 6012
rect 16168 5956 16172 6012
rect 16108 5952 16172 5956
rect 16188 6012 16252 6016
rect 16188 5956 16192 6012
rect 16192 5956 16248 6012
rect 16248 5956 16252 6012
rect 16188 5952 16252 5956
rect 23722 6012 23786 6016
rect 23722 5956 23726 6012
rect 23726 5956 23782 6012
rect 23782 5956 23786 6012
rect 23722 5952 23786 5956
rect 23802 6012 23866 6016
rect 23802 5956 23806 6012
rect 23806 5956 23862 6012
rect 23862 5956 23866 6012
rect 23802 5952 23866 5956
rect 23882 6012 23946 6016
rect 23882 5956 23886 6012
rect 23886 5956 23942 6012
rect 23942 5956 23946 6012
rect 23882 5952 23946 5956
rect 23962 6012 24026 6016
rect 23962 5956 23966 6012
rect 23966 5956 24022 6012
rect 24022 5956 24026 6012
rect 23962 5952 24026 5956
rect 31496 6012 31560 6016
rect 31496 5956 31500 6012
rect 31500 5956 31556 6012
rect 31556 5956 31560 6012
rect 31496 5952 31560 5956
rect 31576 6012 31640 6016
rect 31576 5956 31580 6012
rect 31580 5956 31636 6012
rect 31636 5956 31640 6012
rect 31576 5952 31640 5956
rect 31656 6012 31720 6016
rect 31656 5956 31660 6012
rect 31660 5956 31716 6012
rect 31716 5956 31720 6012
rect 31656 5952 31720 5956
rect 31736 6012 31800 6016
rect 31736 5956 31740 6012
rect 31740 5956 31796 6012
rect 31796 5956 31800 6012
rect 31736 5952 31800 5956
rect 4287 5468 4351 5472
rect 4287 5412 4291 5468
rect 4291 5412 4347 5468
rect 4347 5412 4351 5468
rect 4287 5408 4351 5412
rect 4367 5468 4431 5472
rect 4367 5412 4371 5468
rect 4371 5412 4427 5468
rect 4427 5412 4431 5468
rect 4367 5408 4431 5412
rect 4447 5468 4511 5472
rect 4447 5412 4451 5468
rect 4451 5412 4507 5468
rect 4507 5412 4511 5468
rect 4447 5408 4511 5412
rect 4527 5468 4591 5472
rect 4527 5412 4531 5468
rect 4531 5412 4587 5468
rect 4587 5412 4591 5468
rect 4527 5408 4591 5412
rect 12061 5468 12125 5472
rect 12061 5412 12065 5468
rect 12065 5412 12121 5468
rect 12121 5412 12125 5468
rect 12061 5408 12125 5412
rect 12141 5468 12205 5472
rect 12141 5412 12145 5468
rect 12145 5412 12201 5468
rect 12201 5412 12205 5468
rect 12141 5408 12205 5412
rect 12221 5468 12285 5472
rect 12221 5412 12225 5468
rect 12225 5412 12281 5468
rect 12281 5412 12285 5468
rect 12221 5408 12285 5412
rect 12301 5468 12365 5472
rect 12301 5412 12305 5468
rect 12305 5412 12361 5468
rect 12361 5412 12365 5468
rect 12301 5408 12365 5412
rect 19835 5468 19899 5472
rect 19835 5412 19839 5468
rect 19839 5412 19895 5468
rect 19895 5412 19899 5468
rect 19835 5408 19899 5412
rect 19915 5468 19979 5472
rect 19915 5412 19919 5468
rect 19919 5412 19975 5468
rect 19975 5412 19979 5468
rect 19915 5408 19979 5412
rect 19995 5468 20059 5472
rect 19995 5412 19999 5468
rect 19999 5412 20055 5468
rect 20055 5412 20059 5468
rect 19995 5408 20059 5412
rect 20075 5468 20139 5472
rect 20075 5412 20079 5468
rect 20079 5412 20135 5468
rect 20135 5412 20139 5468
rect 20075 5408 20139 5412
rect 27609 5468 27673 5472
rect 27609 5412 27613 5468
rect 27613 5412 27669 5468
rect 27669 5412 27673 5468
rect 27609 5408 27673 5412
rect 27689 5468 27753 5472
rect 27689 5412 27693 5468
rect 27693 5412 27749 5468
rect 27749 5412 27753 5468
rect 27689 5408 27753 5412
rect 27769 5468 27833 5472
rect 27769 5412 27773 5468
rect 27773 5412 27829 5468
rect 27829 5412 27833 5468
rect 27769 5408 27833 5412
rect 27849 5468 27913 5472
rect 27849 5412 27853 5468
rect 27853 5412 27909 5468
rect 27909 5412 27913 5468
rect 27849 5408 27913 5412
rect 8174 4924 8238 4928
rect 8174 4868 8178 4924
rect 8178 4868 8234 4924
rect 8234 4868 8238 4924
rect 8174 4864 8238 4868
rect 8254 4924 8318 4928
rect 8254 4868 8258 4924
rect 8258 4868 8314 4924
rect 8314 4868 8318 4924
rect 8254 4864 8318 4868
rect 8334 4924 8398 4928
rect 8334 4868 8338 4924
rect 8338 4868 8394 4924
rect 8394 4868 8398 4924
rect 8334 4864 8398 4868
rect 8414 4924 8478 4928
rect 8414 4868 8418 4924
rect 8418 4868 8474 4924
rect 8474 4868 8478 4924
rect 8414 4864 8478 4868
rect 15948 4924 16012 4928
rect 15948 4868 15952 4924
rect 15952 4868 16008 4924
rect 16008 4868 16012 4924
rect 15948 4864 16012 4868
rect 16028 4924 16092 4928
rect 16028 4868 16032 4924
rect 16032 4868 16088 4924
rect 16088 4868 16092 4924
rect 16028 4864 16092 4868
rect 16108 4924 16172 4928
rect 16108 4868 16112 4924
rect 16112 4868 16168 4924
rect 16168 4868 16172 4924
rect 16108 4864 16172 4868
rect 16188 4924 16252 4928
rect 16188 4868 16192 4924
rect 16192 4868 16248 4924
rect 16248 4868 16252 4924
rect 16188 4864 16252 4868
rect 23722 4924 23786 4928
rect 23722 4868 23726 4924
rect 23726 4868 23782 4924
rect 23782 4868 23786 4924
rect 23722 4864 23786 4868
rect 23802 4924 23866 4928
rect 23802 4868 23806 4924
rect 23806 4868 23862 4924
rect 23862 4868 23866 4924
rect 23802 4864 23866 4868
rect 23882 4924 23946 4928
rect 23882 4868 23886 4924
rect 23886 4868 23942 4924
rect 23942 4868 23946 4924
rect 23882 4864 23946 4868
rect 23962 4924 24026 4928
rect 23962 4868 23966 4924
rect 23966 4868 24022 4924
rect 24022 4868 24026 4924
rect 23962 4864 24026 4868
rect 31496 4924 31560 4928
rect 31496 4868 31500 4924
rect 31500 4868 31556 4924
rect 31556 4868 31560 4924
rect 31496 4864 31560 4868
rect 31576 4924 31640 4928
rect 31576 4868 31580 4924
rect 31580 4868 31636 4924
rect 31636 4868 31640 4924
rect 31576 4864 31640 4868
rect 31656 4924 31720 4928
rect 31656 4868 31660 4924
rect 31660 4868 31716 4924
rect 31716 4868 31720 4924
rect 31656 4864 31720 4868
rect 31736 4924 31800 4928
rect 31736 4868 31740 4924
rect 31740 4868 31796 4924
rect 31796 4868 31800 4924
rect 31736 4864 31800 4868
rect 4287 4380 4351 4384
rect 4287 4324 4291 4380
rect 4291 4324 4347 4380
rect 4347 4324 4351 4380
rect 4287 4320 4351 4324
rect 4367 4380 4431 4384
rect 4367 4324 4371 4380
rect 4371 4324 4427 4380
rect 4427 4324 4431 4380
rect 4367 4320 4431 4324
rect 4447 4380 4511 4384
rect 4447 4324 4451 4380
rect 4451 4324 4507 4380
rect 4507 4324 4511 4380
rect 4447 4320 4511 4324
rect 4527 4380 4591 4384
rect 4527 4324 4531 4380
rect 4531 4324 4587 4380
rect 4587 4324 4591 4380
rect 4527 4320 4591 4324
rect 12061 4380 12125 4384
rect 12061 4324 12065 4380
rect 12065 4324 12121 4380
rect 12121 4324 12125 4380
rect 12061 4320 12125 4324
rect 12141 4380 12205 4384
rect 12141 4324 12145 4380
rect 12145 4324 12201 4380
rect 12201 4324 12205 4380
rect 12141 4320 12205 4324
rect 12221 4380 12285 4384
rect 12221 4324 12225 4380
rect 12225 4324 12281 4380
rect 12281 4324 12285 4380
rect 12221 4320 12285 4324
rect 12301 4380 12365 4384
rect 12301 4324 12305 4380
rect 12305 4324 12361 4380
rect 12361 4324 12365 4380
rect 12301 4320 12365 4324
rect 19835 4380 19899 4384
rect 19835 4324 19839 4380
rect 19839 4324 19895 4380
rect 19895 4324 19899 4380
rect 19835 4320 19899 4324
rect 19915 4380 19979 4384
rect 19915 4324 19919 4380
rect 19919 4324 19975 4380
rect 19975 4324 19979 4380
rect 19915 4320 19979 4324
rect 19995 4380 20059 4384
rect 19995 4324 19999 4380
rect 19999 4324 20055 4380
rect 20055 4324 20059 4380
rect 19995 4320 20059 4324
rect 20075 4380 20139 4384
rect 20075 4324 20079 4380
rect 20079 4324 20135 4380
rect 20135 4324 20139 4380
rect 20075 4320 20139 4324
rect 27609 4380 27673 4384
rect 27609 4324 27613 4380
rect 27613 4324 27669 4380
rect 27669 4324 27673 4380
rect 27609 4320 27673 4324
rect 27689 4380 27753 4384
rect 27689 4324 27693 4380
rect 27693 4324 27749 4380
rect 27749 4324 27753 4380
rect 27689 4320 27753 4324
rect 27769 4380 27833 4384
rect 27769 4324 27773 4380
rect 27773 4324 27829 4380
rect 27829 4324 27833 4380
rect 27769 4320 27833 4324
rect 27849 4380 27913 4384
rect 27849 4324 27853 4380
rect 27853 4324 27909 4380
rect 27909 4324 27913 4380
rect 27849 4320 27913 4324
rect 8174 3836 8238 3840
rect 8174 3780 8178 3836
rect 8178 3780 8234 3836
rect 8234 3780 8238 3836
rect 8174 3776 8238 3780
rect 8254 3836 8318 3840
rect 8254 3780 8258 3836
rect 8258 3780 8314 3836
rect 8314 3780 8318 3836
rect 8254 3776 8318 3780
rect 8334 3836 8398 3840
rect 8334 3780 8338 3836
rect 8338 3780 8394 3836
rect 8394 3780 8398 3836
rect 8334 3776 8398 3780
rect 8414 3836 8478 3840
rect 8414 3780 8418 3836
rect 8418 3780 8474 3836
rect 8474 3780 8478 3836
rect 8414 3776 8478 3780
rect 15948 3836 16012 3840
rect 15948 3780 15952 3836
rect 15952 3780 16008 3836
rect 16008 3780 16012 3836
rect 15948 3776 16012 3780
rect 16028 3836 16092 3840
rect 16028 3780 16032 3836
rect 16032 3780 16088 3836
rect 16088 3780 16092 3836
rect 16028 3776 16092 3780
rect 16108 3836 16172 3840
rect 16108 3780 16112 3836
rect 16112 3780 16168 3836
rect 16168 3780 16172 3836
rect 16108 3776 16172 3780
rect 16188 3836 16252 3840
rect 16188 3780 16192 3836
rect 16192 3780 16248 3836
rect 16248 3780 16252 3836
rect 16188 3776 16252 3780
rect 23722 3836 23786 3840
rect 23722 3780 23726 3836
rect 23726 3780 23782 3836
rect 23782 3780 23786 3836
rect 23722 3776 23786 3780
rect 23802 3836 23866 3840
rect 23802 3780 23806 3836
rect 23806 3780 23862 3836
rect 23862 3780 23866 3836
rect 23802 3776 23866 3780
rect 23882 3836 23946 3840
rect 23882 3780 23886 3836
rect 23886 3780 23942 3836
rect 23942 3780 23946 3836
rect 23882 3776 23946 3780
rect 23962 3836 24026 3840
rect 23962 3780 23966 3836
rect 23966 3780 24022 3836
rect 24022 3780 24026 3836
rect 23962 3776 24026 3780
rect 31496 3836 31560 3840
rect 31496 3780 31500 3836
rect 31500 3780 31556 3836
rect 31556 3780 31560 3836
rect 31496 3776 31560 3780
rect 31576 3836 31640 3840
rect 31576 3780 31580 3836
rect 31580 3780 31636 3836
rect 31636 3780 31640 3836
rect 31576 3776 31640 3780
rect 31656 3836 31720 3840
rect 31656 3780 31660 3836
rect 31660 3780 31716 3836
rect 31716 3780 31720 3836
rect 31656 3776 31720 3780
rect 31736 3836 31800 3840
rect 31736 3780 31740 3836
rect 31740 3780 31796 3836
rect 31796 3780 31800 3836
rect 31736 3776 31800 3780
rect 4287 3292 4351 3296
rect 4287 3236 4291 3292
rect 4291 3236 4347 3292
rect 4347 3236 4351 3292
rect 4287 3232 4351 3236
rect 4367 3292 4431 3296
rect 4367 3236 4371 3292
rect 4371 3236 4427 3292
rect 4427 3236 4431 3292
rect 4367 3232 4431 3236
rect 4447 3292 4511 3296
rect 4447 3236 4451 3292
rect 4451 3236 4507 3292
rect 4507 3236 4511 3292
rect 4447 3232 4511 3236
rect 4527 3292 4591 3296
rect 4527 3236 4531 3292
rect 4531 3236 4587 3292
rect 4587 3236 4591 3292
rect 4527 3232 4591 3236
rect 12061 3292 12125 3296
rect 12061 3236 12065 3292
rect 12065 3236 12121 3292
rect 12121 3236 12125 3292
rect 12061 3232 12125 3236
rect 12141 3292 12205 3296
rect 12141 3236 12145 3292
rect 12145 3236 12201 3292
rect 12201 3236 12205 3292
rect 12141 3232 12205 3236
rect 12221 3292 12285 3296
rect 12221 3236 12225 3292
rect 12225 3236 12281 3292
rect 12281 3236 12285 3292
rect 12221 3232 12285 3236
rect 12301 3292 12365 3296
rect 12301 3236 12305 3292
rect 12305 3236 12361 3292
rect 12361 3236 12365 3292
rect 12301 3232 12365 3236
rect 19835 3292 19899 3296
rect 19835 3236 19839 3292
rect 19839 3236 19895 3292
rect 19895 3236 19899 3292
rect 19835 3232 19899 3236
rect 19915 3292 19979 3296
rect 19915 3236 19919 3292
rect 19919 3236 19975 3292
rect 19975 3236 19979 3292
rect 19915 3232 19979 3236
rect 19995 3292 20059 3296
rect 19995 3236 19999 3292
rect 19999 3236 20055 3292
rect 20055 3236 20059 3292
rect 19995 3232 20059 3236
rect 20075 3292 20139 3296
rect 20075 3236 20079 3292
rect 20079 3236 20135 3292
rect 20135 3236 20139 3292
rect 20075 3232 20139 3236
rect 27609 3292 27673 3296
rect 27609 3236 27613 3292
rect 27613 3236 27669 3292
rect 27669 3236 27673 3292
rect 27609 3232 27673 3236
rect 27689 3292 27753 3296
rect 27689 3236 27693 3292
rect 27693 3236 27749 3292
rect 27749 3236 27753 3292
rect 27689 3232 27753 3236
rect 27769 3292 27833 3296
rect 27769 3236 27773 3292
rect 27773 3236 27829 3292
rect 27829 3236 27833 3292
rect 27769 3232 27833 3236
rect 27849 3292 27913 3296
rect 27849 3236 27853 3292
rect 27853 3236 27909 3292
rect 27909 3236 27913 3292
rect 27849 3232 27913 3236
rect 8174 2748 8238 2752
rect 8174 2692 8178 2748
rect 8178 2692 8234 2748
rect 8234 2692 8238 2748
rect 8174 2688 8238 2692
rect 8254 2748 8318 2752
rect 8254 2692 8258 2748
rect 8258 2692 8314 2748
rect 8314 2692 8318 2748
rect 8254 2688 8318 2692
rect 8334 2748 8398 2752
rect 8334 2692 8338 2748
rect 8338 2692 8394 2748
rect 8394 2692 8398 2748
rect 8334 2688 8398 2692
rect 8414 2748 8478 2752
rect 8414 2692 8418 2748
rect 8418 2692 8474 2748
rect 8474 2692 8478 2748
rect 8414 2688 8478 2692
rect 15948 2748 16012 2752
rect 15948 2692 15952 2748
rect 15952 2692 16008 2748
rect 16008 2692 16012 2748
rect 15948 2688 16012 2692
rect 16028 2748 16092 2752
rect 16028 2692 16032 2748
rect 16032 2692 16088 2748
rect 16088 2692 16092 2748
rect 16028 2688 16092 2692
rect 16108 2748 16172 2752
rect 16108 2692 16112 2748
rect 16112 2692 16168 2748
rect 16168 2692 16172 2748
rect 16108 2688 16172 2692
rect 16188 2748 16252 2752
rect 16188 2692 16192 2748
rect 16192 2692 16248 2748
rect 16248 2692 16252 2748
rect 16188 2688 16252 2692
rect 23722 2748 23786 2752
rect 23722 2692 23726 2748
rect 23726 2692 23782 2748
rect 23782 2692 23786 2748
rect 23722 2688 23786 2692
rect 23802 2748 23866 2752
rect 23802 2692 23806 2748
rect 23806 2692 23862 2748
rect 23862 2692 23866 2748
rect 23802 2688 23866 2692
rect 23882 2748 23946 2752
rect 23882 2692 23886 2748
rect 23886 2692 23942 2748
rect 23942 2692 23946 2748
rect 23882 2688 23946 2692
rect 23962 2748 24026 2752
rect 23962 2692 23966 2748
rect 23966 2692 24022 2748
rect 24022 2692 24026 2748
rect 23962 2688 24026 2692
rect 31496 2748 31560 2752
rect 31496 2692 31500 2748
rect 31500 2692 31556 2748
rect 31556 2692 31560 2748
rect 31496 2688 31560 2692
rect 31576 2748 31640 2752
rect 31576 2692 31580 2748
rect 31580 2692 31636 2748
rect 31636 2692 31640 2748
rect 31576 2688 31640 2692
rect 31656 2748 31720 2752
rect 31656 2692 31660 2748
rect 31660 2692 31716 2748
rect 31716 2692 31720 2748
rect 31656 2688 31720 2692
rect 31736 2748 31800 2752
rect 31736 2692 31740 2748
rect 31740 2692 31796 2748
rect 31796 2692 31800 2748
rect 31736 2688 31800 2692
rect 4287 2204 4351 2208
rect 4287 2148 4291 2204
rect 4291 2148 4347 2204
rect 4347 2148 4351 2204
rect 4287 2144 4351 2148
rect 4367 2204 4431 2208
rect 4367 2148 4371 2204
rect 4371 2148 4427 2204
rect 4427 2148 4431 2204
rect 4367 2144 4431 2148
rect 4447 2204 4511 2208
rect 4447 2148 4451 2204
rect 4451 2148 4507 2204
rect 4507 2148 4511 2204
rect 4447 2144 4511 2148
rect 4527 2204 4591 2208
rect 4527 2148 4531 2204
rect 4531 2148 4587 2204
rect 4587 2148 4591 2204
rect 4527 2144 4591 2148
rect 12061 2204 12125 2208
rect 12061 2148 12065 2204
rect 12065 2148 12121 2204
rect 12121 2148 12125 2204
rect 12061 2144 12125 2148
rect 12141 2204 12205 2208
rect 12141 2148 12145 2204
rect 12145 2148 12201 2204
rect 12201 2148 12205 2204
rect 12141 2144 12205 2148
rect 12221 2204 12285 2208
rect 12221 2148 12225 2204
rect 12225 2148 12281 2204
rect 12281 2148 12285 2204
rect 12221 2144 12285 2148
rect 12301 2204 12365 2208
rect 12301 2148 12305 2204
rect 12305 2148 12361 2204
rect 12361 2148 12365 2204
rect 12301 2144 12365 2148
rect 19835 2204 19899 2208
rect 19835 2148 19839 2204
rect 19839 2148 19895 2204
rect 19895 2148 19899 2204
rect 19835 2144 19899 2148
rect 19915 2204 19979 2208
rect 19915 2148 19919 2204
rect 19919 2148 19975 2204
rect 19975 2148 19979 2204
rect 19915 2144 19979 2148
rect 19995 2204 20059 2208
rect 19995 2148 19999 2204
rect 19999 2148 20055 2204
rect 20055 2148 20059 2204
rect 19995 2144 20059 2148
rect 20075 2204 20139 2208
rect 20075 2148 20079 2204
rect 20079 2148 20135 2204
rect 20135 2148 20139 2204
rect 20075 2144 20139 2148
rect 27609 2204 27673 2208
rect 27609 2148 27613 2204
rect 27613 2148 27669 2204
rect 27669 2148 27673 2204
rect 27609 2144 27673 2148
rect 27689 2204 27753 2208
rect 27689 2148 27693 2204
rect 27693 2148 27749 2204
rect 27749 2148 27753 2204
rect 27689 2144 27753 2148
rect 27769 2204 27833 2208
rect 27769 2148 27773 2204
rect 27773 2148 27829 2204
rect 27829 2148 27833 2204
rect 27769 2144 27833 2148
rect 27849 2204 27913 2208
rect 27849 2148 27853 2204
rect 27853 2148 27909 2204
rect 27909 2148 27913 2204
rect 27849 2144 27913 2148
rect 8174 1660 8238 1664
rect 8174 1604 8178 1660
rect 8178 1604 8234 1660
rect 8234 1604 8238 1660
rect 8174 1600 8238 1604
rect 8254 1660 8318 1664
rect 8254 1604 8258 1660
rect 8258 1604 8314 1660
rect 8314 1604 8318 1660
rect 8254 1600 8318 1604
rect 8334 1660 8398 1664
rect 8334 1604 8338 1660
rect 8338 1604 8394 1660
rect 8394 1604 8398 1660
rect 8334 1600 8398 1604
rect 8414 1660 8478 1664
rect 8414 1604 8418 1660
rect 8418 1604 8474 1660
rect 8474 1604 8478 1660
rect 8414 1600 8478 1604
rect 15948 1660 16012 1664
rect 15948 1604 15952 1660
rect 15952 1604 16008 1660
rect 16008 1604 16012 1660
rect 15948 1600 16012 1604
rect 16028 1660 16092 1664
rect 16028 1604 16032 1660
rect 16032 1604 16088 1660
rect 16088 1604 16092 1660
rect 16028 1600 16092 1604
rect 16108 1660 16172 1664
rect 16108 1604 16112 1660
rect 16112 1604 16168 1660
rect 16168 1604 16172 1660
rect 16108 1600 16172 1604
rect 16188 1660 16252 1664
rect 16188 1604 16192 1660
rect 16192 1604 16248 1660
rect 16248 1604 16252 1660
rect 16188 1600 16252 1604
rect 23722 1660 23786 1664
rect 23722 1604 23726 1660
rect 23726 1604 23782 1660
rect 23782 1604 23786 1660
rect 23722 1600 23786 1604
rect 23802 1660 23866 1664
rect 23802 1604 23806 1660
rect 23806 1604 23862 1660
rect 23862 1604 23866 1660
rect 23802 1600 23866 1604
rect 23882 1660 23946 1664
rect 23882 1604 23886 1660
rect 23886 1604 23942 1660
rect 23942 1604 23946 1660
rect 23882 1600 23946 1604
rect 23962 1660 24026 1664
rect 23962 1604 23966 1660
rect 23966 1604 24022 1660
rect 24022 1604 24026 1660
rect 23962 1600 24026 1604
rect 31496 1660 31560 1664
rect 31496 1604 31500 1660
rect 31500 1604 31556 1660
rect 31556 1604 31560 1660
rect 31496 1600 31560 1604
rect 31576 1660 31640 1664
rect 31576 1604 31580 1660
rect 31580 1604 31636 1660
rect 31636 1604 31640 1660
rect 31576 1600 31640 1604
rect 31656 1660 31720 1664
rect 31656 1604 31660 1660
rect 31660 1604 31716 1660
rect 31716 1604 31720 1660
rect 31656 1600 31720 1604
rect 31736 1660 31800 1664
rect 31736 1604 31740 1660
rect 31740 1604 31796 1660
rect 31796 1604 31800 1660
rect 31736 1600 31800 1604
rect 4287 1116 4351 1120
rect 4287 1060 4291 1116
rect 4291 1060 4347 1116
rect 4347 1060 4351 1116
rect 4287 1056 4351 1060
rect 4367 1116 4431 1120
rect 4367 1060 4371 1116
rect 4371 1060 4427 1116
rect 4427 1060 4431 1116
rect 4367 1056 4431 1060
rect 4447 1116 4511 1120
rect 4447 1060 4451 1116
rect 4451 1060 4507 1116
rect 4507 1060 4511 1116
rect 4447 1056 4511 1060
rect 4527 1116 4591 1120
rect 4527 1060 4531 1116
rect 4531 1060 4587 1116
rect 4587 1060 4591 1116
rect 4527 1056 4591 1060
rect 12061 1116 12125 1120
rect 12061 1060 12065 1116
rect 12065 1060 12121 1116
rect 12121 1060 12125 1116
rect 12061 1056 12125 1060
rect 12141 1116 12205 1120
rect 12141 1060 12145 1116
rect 12145 1060 12201 1116
rect 12201 1060 12205 1116
rect 12141 1056 12205 1060
rect 12221 1116 12285 1120
rect 12221 1060 12225 1116
rect 12225 1060 12281 1116
rect 12281 1060 12285 1116
rect 12221 1056 12285 1060
rect 12301 1116 12365 1120
rect 12301 1060 12305 1116
rect 12305 1060 12361 1116
rect 12361 1060 12365 1116
rect 12301 1056 12365 1060
rect 19835 1116 19899 1120
rect 19835 1060 19839 1116
rect 19839 1060 19895 1116
rect 19895 1060 19899 1116
rect 19835 1056 19899 1060
rect 19915 1116 19979 1120
rect 19915 1060 19919 1116
rect 19919 1060 19975 1116
rect 19975 1060 19979 1116
rect 19915 1056 19979 1060
rect 19995 1116 20059 1120
rect 19995 1060 19999 1116
rect 19999 1060 20055 1116
rect 20055 1060 20059 1116
rect 19995 1056 20059 1060
rect 20075 1116 20139 1120
rect 20075 1060 20079 1116
rect 20079 1060 20135 1116
rect 20135 1060 20139 1116
rect 20075 1056 20139 1060
rect 27609 1116 27673 1120
rect 27609 1060 27613 1116
rect 27613 1060 27669 1116
rect 27669 1060 27673 1116
rect 27609 1056 27673 1060
rect 27689 1116 27753 1120
rect 27689 1060 27693 1116
rect 27693 1060 27749 1116
rect 27749 1060 27753 1116
rect 27689 1056 27753 1060
rect 27769 1116 27833 1120
rect 27769 1060 27773 1116
rect 27773 1060 27829 1116
rect 27829 1060 27833 1116
rect 27769 1056 27833 1060
rect 27849 1116 27913 1120
rect 27849 1060 27853 1116
rect 27853 1060 27909 1116
rect 27909 1060 27913 1116
rect 27849 1056 27913 1060
rect 8174 572 8238 576
rect 8174 516 8178 572
rect 8178 516 8234 572
rect 8234 516 8238 572
rect 8174 512 8238 516
rect 8254 572 8318 576
rect 8254 516 8258 572
rect 8258 516 8314 572
rect 8314 516 8318 572
rect 8254 512 8318 516
rect 8334 572 8398 576
rect 8334 516 8338 572
rect 8338 516 8394 572
rect 8394 516 8398 572
rect 8334 512 8398 516
rect 8414 572 8478 576
rect 8414 516 8418 572
rect 8418 516 8474 572
rect 8474 516 8478 572
rect 8414 512 8478 516
rect 15948 572 16012 576
rect 15948 516 15952 572
rect 15952 516 16008 572
rect 16008 516 16012 572
rect 15948 512 16012 516
rect 16028 572 16092 576
rect 16028 516 16032 572
rect 16032 516 16088 572
rect 16088 516 16092 572
rect 16028 512 16092 516
rect 16108 572 16172 576
rect 16108 516 16112 572
rect 16112 516 16168 572
rect 16168 516 16172 572
rect 16108 512 16172 516
rect 16188 572 16252 576
rect 16188 516 16192 572
rect 16192 516 16248 572
rect 16248 516 16252 572
rect 16188 512 16252 516
rect 23722 572 23786 576
rect 23722 516 23726 572
rect 23726 516 23782 572
rect 23782 516 23786 572
rect 23722 512 23786 516
rect 23802 572 23866 576
rect 23802 516 23806 572
rect 23806 516 23862 572
rect 23862 516 23866 572
rect 23802 512 23866 516
rect 23882 572 23946 576
rect 23882 516 23886 572
rect 23886 516 23942 572
rect 23942 516 23946 572
rect 23882 512 23946 516
rect 23962 572 24026 576
rect 23962 516 23966 572
rect 23966 516 24022 572
rect 24022 516 24026 572
rect 23962 512 24026 516
rect 31496 572 31560 576
rect 31496 516 31500 572
rect 31500 516 31556 572
rect 31556 516 31560 572
rect 31496 512 31560 516
rect 31576 572 31640 576
rect 31576 516 31580 572
rect 31580 516 31636 572
rect 31636 516 31640 572
rect 31576 512 31640 516
rect 31656 572 31720 576
rect 31656 516 31660 572
rect 31660 516 31716 572
rect 31716 516 31720 572
rect 31656 512 31720 516
rect 31736 572 31800 576
rect 31736 516 31740 572
rect 31740 516 31796 572
rect 31796 516 31800 572
rect 31736 512 31800 516
<< metal4 >>
rect 798 21861 858 22304
rect 1534 21861 1594 22304
rect 2270 21861 2330 22304
rect 3006 21861 3066 22304
rect 3742 21861 3802 22304
rect 4478 21997 4538 22304
rect 4475 21996 4541 21997
rect 4475 21932 4476 21996
rect 4540 21932 4541 21996
rect 4475 21931 4541 21932
rect 5214 21861 5274 22304
rect 5950 21861 6010 22304
rect 6686 21861 6746 22304
rect 7422 21861 7482 22304
rect 8158 21997 8218 22304
rect 8155 21996 8221 21997
rect 8155 21932 8156 21996
rect 8220 21932 8221 21996
rect 8155 21931 8221 21932
rect 8894 21861 8954 22304
rect 9630 21861 9690 22304
rect 10366 21861 10426 22304
rect 11102 21861 11162 22304
rect 11838 21861 11898 22304
rect 12574 21861 12634 22304
rect 13310 21861 13370 22304
rect 14046 21861 14106 22304
rect 14782 21861 14842 22304
rect 15518 21861 15578 22304
rect 16254 21997 16314 22304
rect 16251 21996 16317 21997
rect 16251 21932 16252 21996
rect 16316 21932 16317 21996
rect 16251 21931 16317 21932
rect 16990 21861 17050 22304
rect 795 21860 861 21861
rect 795 21796 796 21860
rect 860 21796 861 21860
rect 795 21795 861 21796
rect 1531 21860 1597 21861
rect 1531 21796 1532 21860
rect 1596 21796 1597 21860
rect 1531 21795 1597 21796
rect 2267 21860 2333 21861
rect 2267 21796 2268 21860
rect 2332 21796 2333 21860
rect 2267 21795 2333 21796
rect 3003 21860 3069 21861
rect 3003 21796 3004 21860
rect 3068 21796 3069 21860
rect 3003 21795 3069 21796
rect 3739 21860 3805 21861
rect 3739 21796 3740 21860
rect 3804 21796 3805 21860
rect 5211 21860 5277 21861
rect 3739 21795 3805 21796
rect 4279 21792 4599 21808
rect 5211 21796 5212 21860
rect 5276 21796 5277 21860
rect 5211 21795 5277 21796
rect 5947 21860 6013 21861
rect 5947 21796 5948 21860
rect 6012 21796 6013 21860
rect 5947 21795 6013 21796
rect 6683 21860 6749 21861
rect 6683 21796 6684 21860
rect 6748 21796 6749 21860
rect 6683 21795 6749 21796
rect 7419 21860 7485 21861
rect 7419 21796 7420 21860
rect 7484 21796 7485 21860
rect 8891 21860 8957 21861
rect 7419 21795 7485 21796
rect 4279 21728 4287 21792
rect 4351 21728 4367 21792
rect 4431 21728 4447 21792
rect 4511 21728 4527 21792
rect 4591 21728 4599 21792
rect 4279 20704 4599 21728
rect 4279 20640 4287 20704
rect 4351 20640 4367 20704
rect 4431 20640 4447 20704
rect 4511 20640 4527 20704
rect 4591 20640 4599 20704
rect 4279 19616 4599 20640
rect 4279 19552 4287 19616
rect 4351 19552 4367 19616
rect 4431 19552 4447 19616
rect 4511 19552 4527 19616
rect 4591 19552 4599 19616
rect 4279 18528 4599 19552
rect 4279 18464 4287 18528
rect 4351 18464 4367 18528
rect 4431 18464 4447 18528
rect 4511 18464 4527 18528
rect 4591 18464 4599 18528
rect 4279 17440 4599 18464
rect 4279 17376 4287 17440
rect 4351 17376 4367 17440
rect 4431 17376 4447 17440
rect 4511 17376 4527 17440
rect 4591 17376 4599 17440
rect 4279 16352 4599 17376
rect 4279 16288 4287 16352
rect 4351 16288 4367 16352
rect 4431 16288 4447 16352
rect 4511 16288 4527 16352
rect 4591 16288 4599 16352
rect 4279 15264 4599 16288
rect 4279 15200 4287 15264
rect 4351 15200 4367 15264
rect 4431 15200 4447 15264
rect 4511 15200 4527 15264
rect 4591 15200 4599 15264
rect 4279 14176 4599 15200
rect 4279 14112 4287 14176
rect 4351 14112 4367 14176
rect 4431 14112 4447 14176
rect 4511 14112 4527 14176
rect 4591 14112 4599 14176
rect 4279 13088 4599 14112
rect 4279 13024 4287 13088
rect 4351 13024 4367 13088
rect 4431 13024 4447 13088
rect 4511 13024 4527 13088
rect 4591 13024 4599 13088
rect 4279 12000 4599 13024
rect 4279 11936 4287 12000
rect 4351 11936 4367 12000
rect 4431 11936 4447 12000
rect 4511 11936 4527 12000
rect 4591 11936 4599 12000
rect 4279 10912 4599 11936
rect 4279 10848 4287 10912
rect 4351 10848 4367 10912
rect 4431 10848 4447 10912
rect 4511 10848 4527 10912
rect 4591 10848 4599 10912
rect 4279 9824 4599 10848
rect 4279 9760 4287 9824
rect 4351 9760 4367 9824
rect 4431 9760 4447 9824
rect 4511 9760 4527 9824
rect 4591 9760 4599 9824
rect 4279 8736 4599 9760
rect 4279 8672 4287 8736
rect 4351 8672 4367 8736
rect 4431 8672 4447 8736
rect 4511 8672 4527 8736
rect 4591 8672 4599 8736
rect 4279 7648 4599 8672
rect 4279 7584 4287 7648
rect 4351 7584 4367 7648
rect 4431 7584 4447 7648
rect 4511 7584 4527 7648
rect 4591 7584 4599 7648
rect 4279 6560 4599 7584
rect 4279 6496 4287 6560
rect 4351 6496 4367 6560
rect 4431 6496 4447 6560
rect 4511 6496 4527 6560
rect 4591 6496 4599 6560
rect 4279 5472 4599 6496
rect 4279 5408 4287 5472
rect 4351 5408 4367 5472
rect 4431 5408 4447 5472
rect 4511 5408 4527 5472
rect 4591 5408 4599 5472
rect 4279 4384 4599 5408
rect 4279 4320 4287 4384
rect 4351 4320 4367 4384
rect 4431 4320 4447 4384
rect 4511 4320 4527 4384
rect 4591 4320 4599 4384
rect 4279 3296 4599 4320
rect 4279 3232 4287 3296
rect 4351 3232 4367 3296
rect 4431 3232 4447 3296
rect 4511 3232 4527 3296
rect 4591 3232 4599 3296
rect 4279 2208 4599 3232
rect 4279 2144 4287 2208
rect 4351 2144 4367 2208
rect 4431 2144 4447 2208
rect 4511 2144 4527 2208
rect 4591 2144 4599 2208
rect 4279 1120 4599 2144
rect 4279 1056 4287 1120
rect 4351 1056 4367 1120
rect 4431 1056 4447 1120
rect 4511 1056 4527 1120
rect 4591 1056 4599 1120
rect 4279 496 4599 1056
rect 8166 21248 8486 21808
rect 8891 21796 8892 21860
rect 8956 21796 8957 21860
rect 8891 21795 8957 21796
rect 9627 21860 9693 21861
rect 9627 21796 9628 21860
rect 9692 21796 9693 21860
rect 9627 21795 9693 21796
rect 10363 21860 10429 21861
rect 10363 21796 10364 21860
rect 10428 21796 10429 21860
rect 10363 21795 10429 21796
rect 11099 21860 11165 21861
rect 11099 21796 11100 21860
rect 11164 21796 11165 21860
rect 11099 21795 11165 21796
rect 11835 21860 11901 21861
rect 11835 21796 11836 21860
rect 11900 21796 11901 21860
rect 12571 21860 12637 21861
rect 11835 21795 11901 21796
rect 8166 21184 8174 21248
rect 8238 21184 8254 21248
rect 8318 21184 8334 21248
rect 8398 21184 8414 21248
rect 8478 21184 8486 21248
rect 8166 20160 8486 21184
rect 8166 20096 8174 20160
rect 8238 20096 8254 20160
rect 8318 20096 8334 20160
rect 8398 20096 8414 20160
rect 8478 20096 8486 20160
rect 8166 19072 8486 20096
rect 8166 19008 8174 19072
rect 8238 19008 8254 19072
rect 8318 19008 8334 19072
rect 8398 19008 8414 19072
rect 8478 19008 8486 19072
rect 8166 17984 8486 19008
rect 8166 17920 8174 17984
rect 8238 17920 8254 17984
rect 8318 17920 8334 17984
rect 8398 17920 8414 17984
rect 8478 17920 8486 17984
rect 8166 16896 8486 17920
rect 8166 16832 8174 16896
rect 8238 16832 8254 16896
rect 8318 16832 8334 16896
rect 8398 16832 8414 16896
rect 8478 16832 8486 16896
rect 8166 15808 8486 16832
rect 8166 15744 8174 15808
rect 8238 15744 8254 15808
rect 8318 15744 8334 15808
rect 8398 15744 8414 15808
rect 8478 15744 8486 15808
rect 8166 14720 8486 15744
rect 8166 14656 8174 14720
rect 8238 14656 8254 14720
rect 8318 14656 8334 14720
rect 8398 14656 8414 14720
rect 8478 14656 8486 14720
rect 8166 13632 8486 14656
rect 8166 13568 8174 13632
rect 8238 13568 8254 13632
rect 8318 13568 8334 13632
rect 8398 13568 8414 13632
rect 8478 13568 8486 13632
rect 8166 12544 8486 13568
rect 8166 12480 8174 12544
rect 8238 12480 8254 12544
rect 8318 12480 8334 12544
rect 8398 12480 8414 12544
rect 8478 12480 8486 12544
rect 8166 11456 8486 12480
rect 8166 11392 8174 11456
rect 8238 11392 8254 11456
rect 8318 11392 8334 11456
rect 8398 11392 8414 11456
rect 8478 11392 8486 11456
rect 8166 10368 8486 11392
rect 8166 10304 8174 10368
rect 8238 10304 8254 10368
rect 8318 10304 8334 10368
rect 8398 10304 8414 10368
rect 8478 10304 8486 10368
rect 8166 9280 8486 10304
rect 8166 9216 8174 9280
rect 8238 9216 8254 9280
rect 8318 9216 8334 9280
rect 8398 9216 8414 9280
rect 8478 9216 8486 9280
rect 8166 8192 8486 9216
rect 8166 8128 8174 8192
rect 8238 8128 8254 8192
rect 8318 8128 8334 8192
rect 8398 8128 8414 8192
rect 8478 8128 8486 8192
rect 8166 7104 8486 8128
rect 8166 7040 8174 7104
rect 8238 7040 8254 7104
rect 8318 7040 8334 7104
rect 8398 7040 8414 7104
rect 8478 7040 8486 7104
rect 8166 6016 8486 7040
rect 8166 5952 8174 6016
rect 8238 5952 8254 6016
rect 8318 5952 8334 6016
rect 8398 5952 8414 6016
rect 8478 5952 8486 6016
rect 8166 4928 8486 5952
rect 8166 4864 8174 4928
rect 8238 4864 8254 4928
rect 8318 4864 8334 4928
rect 8398 4864 8414 4928
rect 8478 4864 8486 4928
rect 8166 3840 8486 4864
rect 8166 3776 8174 3840
rect 8238 3776 8254 3840
rect 8318 3776 8334 3840
rect 8398 3776 8414 3840
rect 8478 3776 8486 3840
rect 8166 2752 8486 3776
rect 8166 2688 8174 2752
rect 8238 2688 8254 2752
rect 8318 2688 8334 2752
rect 8398 2688 8414 2752
rect 8478 2688 8486 2752
rect 8166 1664 8486 2688
rect 8166 1600 8174 1664
rect 8238 1600 8254 1664
rect 8318 1600 8334 1664
rect 8398 1600 8414 1664
rect 8478 1600 8486 1664
rect 8166 576 8486 1600
rect 8166 512 8174 576
rect 8238 512 8254 576
rect 8318 512 8334 576
rect 8398 512 8414 576
rect 8478 512 8486 576
rect 8166 496 8486 512
rect 12053 21792 12373 21808
rect 12571 21796 12572 21860
rect 12636 21796 12637 21860
rect 12571 21795 12637 21796
rect 13307 21860 13373 21861
rect 13307 21796 13308 21860
rect 13372 21796 13373 21860
rect 13307 21795 13373 21796
rect 14043 21860 14109 21861
rect 14043 21796 14044 21860
rect 14108 21796 14109 21860
rect 14043 21795 14109 21796
rect 14779 21860 14845 21861
rect 14779 21796 14780 21860
rect 14844 21796 14845 21860
rect 14779 21795 14845 21796
rect 15515 21860 15581 21861
rect 15515 21796 15516 21860
rect 15580 21796 15581 21860
rect 16987 21860 17053 21861
rect 15515 21795 15581 21796
rect 12053 21728 12061 21792
rect 12125 21728 12141 21792
rect 12205 21728 12221 21792
rect 12285 21728 12301 21792
rect 12365 21728 12373 21792
rect 12053 20704 12373 21728
rect 12053 20640 12061 20704
rect 12125 20640 12141 20704
rect 12205 20640 12221 20704
rect 12285 20640 12301 20704
rect 12365 20640 12373 20704
rect 12053 19616 12373 20640
rect 12053 19552 12061 19616
rect 12125 19552 12141 19616
rect 12205 19552 12221 19616
rect 12285 19552 12301 19616
rect 12365 19552 12373 19616
rect 12053 18528 12373 19552
rect 12053 18464 12061 18528
rect 12125 18464 12141 18528
rect 12205 18464 12221 18528
rect 12285 18464 12301 18528
rect 12365 18464 12373 18528
rect 12053 17440 12373 18464
rect 12053 17376 12061 17440
rect 12125 17376 12141 17440
rect 12205 17376 12221 17440
rect 12285 17376 12301 17440
rect 12365 17376 12373 17440
rect 12053 16352 12373 17376
rect 12053 16288 12061 16352
rect 12125 16288 12141 16352
rect 12205 16288 12221 16352
rect 12285 16288 12301 16352
rect 12365 16288 12373 16352
rect 12053 15264 12373 16288
rect 12053 15200 12061 15264
rect 12125 15200 12141 15264
rect 12205 15200 12221 15264
rect 12285 15200 12301 15264
rect 12365 15200 12373 15264
rect 12053 14176 12373 15200
rect 12053 14112 12061 14176
rect 12125 14112 12141 14176
rect 12205 14112 12221 14176
rect 12285 14112 12301 14176
rect 12365 14112 12373 14176
rect 12053 13088 12373 14112
rect 12053 13024 12061 13088
rect 12125 13024 12141 13088
rect 12205 13024 12221 13088
rect 12285 13024 12301 13088
rect 12365 13024 12373 13088
rect 12053 12000 12373 13024
rect 12053 11936 12061 12000
rect 12125 11936 12141 12000
rect 12205 11936 12221 12000
rect 12285 11936 12301 12000
rect 12365 11936 12373 12000
rect 12053 10912 12373 11936
rect 12053 10848 12061 10912
rect 12125 10848 12141 10912
rect 12205 10848 12221 10912
rect 12285 10848 12301 10912
rect 12365 10848 12373 10912
rect 12053 9824 12373 10848
rect 12053 9760 12061 9824
rect 12125 9760 12141 9824
rect 12205 9760 12221 9824
rect 12285 9760 12301 9824
rect 12365 9760 12373 9824
rect 12053 8736 12373 9760
rect 12053 8672 12061 8736
rect 12125 8672 12141 8736
rect 12205 8672 12221 8736
rect 12285 8672 12301 8736
rect 12365 8672 12373 8736
rect 12053 7648 12373 8672
rect 12053 7584 12061 7648
rect 12125 7584 12141 7648
rect 12205 7584 12221 7648
rect 12285 7584 12301 7648
rect 12365 7584 12373 7648
rect 12053 6560 12373 7584
rect 12053 6496 12061 6560
rect 12125 6496 12141 6560
rect 12205 6496 12221 6560
rect 12285 6496 12301 6560
rect 12365 6496 12373 6560
rect 12053 5472 12373 6496
rect 12053 5408 12061 5472
rect 12125 5408 12141 5472
rect 12205 5408 12221 5472
rect 12285 5408 12301 5472
rect 12365 5408 12373 5472
rect 12053 4384 12373 5408
rect 12053 4320 12061 4384
rect 12125 4320 12141 4384
rect 12205 4320 12221 4384
rect 12285 4320 12301 4384
rect 12365 4320 12373 4384
rect 12053 3296 12373 4320
rect 12053 3232 12061 3296
rect 12125 3232 12141 3296
rect 12205 3232 12221 3296
rect 12285 3232 12301 3296
rect 12365 3232 12373 3296
rect 12053 2208 12373 3232
rect 12053 2144 12061 2208
rect 12125 2144 12141 2208
rect 12205 2144 12221 2208
rect 12285 2144 12301 2208
rect 12365 2144 12373 2208
rect 12053 1120 12373 2144
rect 12053 1056 12061 1120
rect 12125 1056 12141 1120
rect 12205 1056 12221 1120
rect 12285 1056 12301 1120
rect 12365 1056 12373 1120
rect 12053 496 12373 1056
rect 15940 21248 16260 21808
rect 16987 21796 16988 21860
rect 17052 21796 17053 21860
rect 16987 21795 17053 21796
rect 15940 21184 15948 21248
rect 16012 21184 16028 21248
rect 16092 21184 16108 21248
rect 16172 21184 16188 21248
rect 16252 21184 16260 21248
rect 15940 20160 16260 21184
rect 15940 20096 15948 20160
rect 16012 20096 16028 20160
rect 16092 20096 16108 20160
rect 16172 20096 16188 20160
rect 16252 20096 16260 20160
rect 15940 19072 16260 20096
rect 17726 19277 17786 22304
rect 18462 22104 18522 22304
rect 19198 22104 19258 22304
rect 19934 22104 19994 22304
rect 20670 22104 20730 22304
rect 21406 22104 21466 22304
rect 22142 22104 22202 22304
rect 22878 22104 22938 22304
rect 23614 22104 23674 22304
rect 24350 22104 24410 22304
rect 25086 22104 25146 22304
rect 25822 22104 25882 22304
rect 26558 22104 26618 22304
rect 27294 22104 27354 22304
rect 28030 22104 28090 22304
rect 28766 22130 28826 22304
rect 28947 22268 29013 22269
rect 28947 22204 28948 22268
rect 29012 22204 29013 22268
rect 28947 22203 29013 22204
rect 28950 22130 29010 22203
rect 28766 22070 29010 22130
rect 29502 21861 29562 22304
rect 30238 22104 30298 22304
rect 30974 22104 31034 22304
rect 31710 22104 31770 22304
rect 29499 21860 29565 21861
rect 19827 21792 20147 21808
rect 19827 21728 19835 21792
rect 19899 21728 19915 21792
rect 19979 21728 19995 21792
rect 20059 21728 20075 21792
rect 20139 21728 20147 21792
rect 19827 20704 20147 21728
rect 19827 20640 19835 20704
rect 19899 20640 19915 20704
rect 19979 20640 19995 20704
rect 20059 20640 20075 20704
rect 20139 20640 20147 20704
rect 19827 19616 20147 20640
rect 19827 19552 19835 19616
rect 19899 19552 19915 19616
rect 19979 19552 19995 19616
rect 20059 19552 20075 19616
rect 20139 19552 20147 19616
rect 17723 19276 17789 19277
rect 17723 19212 17724 19276
rect 17788 19212 17789 19276
rect 17723 19211 17789 19212
rect 15940 19008 15948 19072
rect 16012 19008 16028 19072
rect 16092 19008 16108 19072
rect 16172 19008 16188 19072
rect 16252 19008 16260 19072
rect 15940 17984 16260 19008
rect 15940 17920 15948 17984
rect 16012 17920 16028 17984
rect 16092 17920 16108 17984
rect 16172 17920 16188 17984
rect 16252 17920 16260 17984
rect 15940 16896 16260 17920
rect 15940 16832 15948 16896
rect 16012 16832 16028 16896
rect 16092 16832 16108 16896
rect 16172 16832 16188 16896
rect 16252 16832 16260 16896
rect 15940 15808 16260 16832
rect 15940 15744 15948 15808
rect 16012 15744 16028 15808
rect 16092 15744 16108 15808
rect 16172 15744 16188 15808
rect 16252 15744 16260 15808
rect 15940 14720 16260 15744
rect 15940 14656 15948 14720
rect 16012 14656 16028 14720
rect 16092 14656 16108 14720
rect 16172 14656 16188 14720
rect 16252 14656 16260 14720
rect 15940 13632 16260 14656
rect 15940 13568 15948 13632
rect 16012 13568 16028 13632
rect 16092 13568 16108 13632
rect 16172 13568 16188 13632
rect 16252 13568 16260 13632
rect 15940 12544 16260 13568
rect 15940 12480 15948 12544
rect 16012 12480 16028 12544
rect 16092 12480 16108 12544
rect 16172 12480 16188 12544
rect 16252 12480 16260 12544
rect 15940 11456 16260 12480
rect 15940 11392 15948 11456
rect 16012 11392 16028 11456
rect 16092 11392 16108 11456
rect 16172 11392 16188 11456
rect 16252 11392 16260 11456
rect 15940 10368 16260 11392
rect 15940 10304 15948 10368
rect 16012 10304 16028 10368
rect 16092 10304 16108 10368
rect 16172 10304 16188 10368
rect 16252 10304 16260 10368
rect 15940 9280 16260 10304
rect 15940 9216 15948 9280
rect 16012 9216 16028 9280
rect 16092 9216 16108 9280
rect 16172 9216 16188 9280
rect 16252 9216 16260 9280
rect 15940 8192 16260 9216
rect 15940 8128 15948 8192
rect 16012 8128 16028 8192
rect 16092 8128 16108 8192
rect 16172 8128 16188 8192
rect 16252 8128 16260 8192
rect 15940 7104 16260 8128
rect 15940 7040 15948 7104
rect 16012 7040 16028 7104
rect 16092 7040 16108 7104
rect 16172 7040 16188 7104
rect 16252 7040 16260 7104
rect 15940 6016 16260 7040
rect 15940 5952 15948 6016
rect 16012 5952 16028 6016
rect 16092 5952 16108 6016
rect 16172 5952 16188 6016
rect 16252 5952 16260 6016
rect 15940 4928 16260 5952
rect 15940 4864 15948 4928
rect 16012 4864 16028 4928
rect 16092 4864 16108 4928
rect 16172 4864 16188 4928
rect 16252 4864 16260 4928
rect 15940 3840 16260 4864
rect 15940 3776 15948 3840
rect 16012 3776 16028 3840
rect 16092 3776 16108 3840
rect 16172 3776 16188 3840
rect 16252 3776 16260 3840
rect 15940 2752 16260 3776
rect 15940 2688 15948 2752
rect 16012 2688 16028 2752
rect 16092 2688 16108 2752
rect 16172 2688 16188 2752
rect 16252 2688 16260 2752
rect 15940 1664 16260 2688
rect 15940 1600 15948 1664
rect 16012 1600 16028 1664
rect 16092 1600 16108 1664
rect 16172 1600 16188 1664
rect 16252 1600 16260 1664
rect 15940 576 16260 1600
rect 15940 512 15948 576
rect 16012 512 16028 576
rect 16092 512 16108 576
rect 16172 512 16188 576
rect 16252 512 16260 576
rect 15940 496 16260 512
rect 19827 18528 20147 19552
rect 19827 18464 19835 18528
rect 19899 18464 19915 18528
rect 19979 18464 19995 18528
rect 20059 18464 20075 18528
rect 20139 18464 20147 18528
rect 19827 17440 20147 18464
rect 19827 17376 19835 17440
rect 19899 17376 19915 17440
rect 19979 17376 19995 17440
rect 20059 17376 20075 17440
rect 20139 17376 20147 17440
rect 19827 16352 20147 17376
rect 19827 16288 19835 16352
rect 19899 16288 19915 16352
rect 19979 16288 19995 16352
rect 20059 16288 20075 16352
rect 20139 16288 20147 16352
rect 19827 15264 20147 16288
rect 19827 15200 19835 15264
rect 19899 15200 19915 15264
rect 19979 15200 19995 15264
rect 20059 15200 20075 15264
rect 20139 15200 20147 15264
rect 19827 14176 20147 15200
rect 19827 14112 19835 14176
rect 19899 14112 19915 14176
rect 19979 14112 19995 14176
rect 20059 14112 20075 14176
rect 20139 14112 20147 14176
rect 19827 13088 20147 14112
rect 19827 13024 19835 13088
rect 19899 13024 19915 13088
rect 19979 13024 19995 13088
rect 20059 13024 20075 13088
rect 20139 13024 20147 13088
rect 19827 12000 20147 13024
rect 19827 11936 19835 12000
rect 19899 11936 19915 12000
rect 19979 11936 19995 12000
rect 20059 11936 20075 12000
rect 20139 11936 20147 12000
rect 19827 10912 20147 11936
rect 19827 10848 19835 10912
rect 19899 10848 19915 10912
rect 19979 10848 19995 10912
rect 20059 10848 20075 10912
rect 20139 10848 20147 10912
rect 19827 9824 20147 10848
rect 19827 9760 19835 9824
rect 19899 9760 19915 9824
rect 19979 9760 19995 9824
rect 20059 9760 20075 9824
rect 20139 9760 20147 9824
rect 19827 8736 20147 9760
rect 19827 8672 19835 8736
rect 19899 8672 19915 8736
rect 19979 8672 19995 8736
rect 20059 8672 20075 8736
rect 20139 8672 20147 8736
rect 19827 7648 20147 8672
rect 19827 7584 19835 7648
rect 19899 7584 19915 7648
rect 19979 7584 19995 7648
rect 20059 7584 20075 7648
rect 20139 7584 20147 7648
rect 19827 6560 20147 7584
rect 19827 6496 19835 6560
rect 19899 6496 19915 6560
rect 19979 6496 19995 6560
rect 20059 6496 20075 6560
rect 20139 6496 20147 6560
rect 19827 5472 20147 6496
rect 19827 5408 19835 5472
rect 19899 5408 19915 5472
rect 19979 5408 19995 5472
rect 20059 5408 20075 5472
rect 20139 5408 20147 5472
rect 19827 4384 20147 5408
rect 19827 4320 19835 4384
rect 19899 4320 19915 4384
rect 19979 4320 19995 4384
rect 20059 4320 20075 4384
rect 20139 4320 20147 4384
rect 19827 3296 20147 4320
rect 19827 3232 19835 3296
rect 19899 3232 19915 3296
rect 19979 3232 19995 3296
rect 20059 3232 20075 3296
rect 20139 3232 20147 3296
rect 19827 2208 20147 3232
rect 19827 2144 19835 2208
rect 19899 2144 19915 2208
rect 19979 2144 19995 2208
rect 20059 2144 20075 2208
rect 20139 2144 20147 2208
rect 19827 1120 20147 2144
rect 19827 1056 19835 1120
rect 19899 1056 19915 1120
rect 19979 1056 19995 1120
rect 20059 1056 20075 1120
rect 20139 1056 20147 1120
rect 19827 496 20147 1056
rect 23714 21248 24034 21808
rect 23714 21184 23722 21248
rect 23786 21184 23802 21248
rect 23866 21184 23882 21248
rect 23946 21184 23962 21248
rect 24026 21184 24034 21248
rect 23714 20160 24034 21184
rect 23714 20096 23722 20160
rect 23786 20096 23802 20160
rect 23866 20096 23882 20160
rect 23946 20096 23962 20160
rect 24026 20096 24034 20160
rect 23714 19072 24034 20096
rect 23714 19008 23722 19072
rect 23786 19008 23802 19072
rect 23866 19008 23882 19072
rect 23946 19008 23962 19072
rect 24026 19008 24034 19072
rect 23714 17984 24034 19008
rect 23714 17920 23722 17984
rect 23786 17920 23802 17984
rect 23866 17920 23882 17984
rect 23946 17920 23962 17984
rect 24026 17920 24034 17984
rect 23714 16896 24034 17920
rect 23714 16832 23722 16896
rect 23786 16832 23802 16896
rect 23866 16832 23882 16896
rect 23946 16832 23962 16896
rect 24026 16832 24034 16896
rect 23714 15808 24034 16832
rect 23714 15744 23722 15808
rect 23786 15744 23802 15808
rect 23866 15744 23882 15808
rect 23946 15744 23962 15808
rect 24026 15744 24034 15808
rect 23714 14720 24034 15744
rect 23714 14656 23722 14720
rect 23786 14656 23802 14720
rect 23866 14656 23882 14720
rect 23946 14656 23962 14720
rect 24026 14656 24034 14720
rect 23714 13632 24034 14656
rect 23714 13568 23722 13632
rect 23786 13568 23802 13632
rect 23866 13568 23882 13632
rect 23946 13568 23962 13632
rect 24026 13568 24034 13632
rect 23714 12544 24034 13568
rect 23714 12480 23722 12544
rect 23786 12480 23802 12544
rect 23866 12480 23882 12544
rect 23946 12480 23962 12544
rect 24026 12480 24034 12544
rect 23714 11456 24034 12480
rect 23714 11392 23722 11456
rect 23786 11392 23802 11456
rect 23866 11392 23882 11456
rect 23946 11392 23962 11456
rect 24026 11392 24034 11456
rect 23714 10368 24034 11392
rect 23714 10304 23722 10368
rect 23786 10304 23802 10368
rect 23866 10304 23882 10368
rect 23946 10304 23962 10368
rect 24026 10304 24034 10368
rect 23714 9280 24034 10304
rect 23714 9216 23722 9280
rect 23786 9216 23802 9280
rect 23866 9216 23882 9280
rect 23946 9216 23962 9280
rect 24026 9216 24034 9280
rect 23714 8192 24034 9216
rect 23714 8128 23722 8192
rect 23786 8128 23802 8192
rect 23866 8128 23882 8192
rect 23946 8128 23962 8192
rect 24026 8128 24034 8192
rect 23714 7104 24034 8128
rect 23714 7040 23722 7104
rect 23786 7040 23802 7104
rect 23866 7040 23882 7104
rect 23946 7040 23962 7104
rect 24026 7040 24034 7104
rect 23714 6016 24034 7040
rect 23714 5952 23722 6016
rect 23786 5952 23802 6016
rect 23866 5952 23882 6016
rect 23946 5952 23962 6016
rect 24026 5952 24034 6016
rect 23714 4928 24034 5952
rect 23714 4864 23722 4928
rect 23786 4864 23802 4928
rect 23866 4864 23882 4928
rect 23946 4864 23962 4928
rect 24026 4864 24034 4928
rect 23714 3840 24034 4864
rect 23714 3776 23722 3840
rect 23786 3776 23802 3840
rect 23866 3776 23882 3840
rect 23946 3776 23962 3840
rect 24026 3776 24034 3840
rect 23714 2752 24034 3776
rect 23714 2688 23722 2752
rect 23786 2688 23802 2752
rect 23866 2688 23882 2752
rect 23946 2688 23962 2752
rect 24026 2688 24034 2752
rect 23714 1664 24034 2688
rect 23714 1600 23722 1664
rect 23786 1600 23802 1664
rect 23866 1600 23882 1664
rect 23946 1600 23962 1664
rect 24026 1600 24034 1664
rect 23714 576 24034 1600
rect 23714 512 23722 576
rect 23786 512 23802 576
rect 23866 512 23882 576
rect 23946 512 23962 576
rect 24026 512 24034 576
rect 23714 496 24034 512
rect 27601 21792 27921 21808
rect 29499 21796 29500 21860
rect 29564 21796 29565 21860
rect 29499 21795 29565 21796
rect 27601 21728 27609 21792
rect 27673 21728 27689 21792
rect 27753 21728 27769 21792
rect 27833 21728 27849 21792
rect 27913 21728 27921 21792
rect 27601 20704 27921 21728
rect 27601 20640 27609 20704
rect 27673 20640 27689 20704
rect 27753 20640 27769 20704
rect 27833 20640 27849 20704
rect 27913 20640 27921 20704
rect 27601 19616 27921 20640
rect 27601 19552 27609 19616
rect 27673 19552 27689 19616
rect 27753 19552 27769 19616
rect 27833 19552 27849 19616
rect 27913 19552 27921 19616
rect 27601 18528 27921 19552
rect 27601 18464 27609 18528
rect 27673 18464 27689 18528
rect 27753 18464 27769 18528
rect 27833 18464 27849 18528
rect 27913 18464 27921 18528
rect 27601 17440 27921 18464
rect 27601 17376 27609 17440
rect 27673 17376 27689 17440
rect 27753 17376 27769 17440
rect 27833 17376 27849 17440
rect 27913 17376 27921 17440
rect 27601 16352 27921 17376
rect 27601 16288 27609 16352
rect 27673 16288 27689 16352
rect 27753 16288 27769 16352
rect 27833 16288 27849 16352
rect 27913 16288 27921 16352
rect 27601 15264 27921 16288
rect 27601 15200 27609 15264
rect 27673 15200 27689 15264
rect 27753 15200 27769 15264
rect 27833 15200 27849 15264
rect 27913 15200 27921 15264
rect 27601 14176 27921 15200
rect 27601 14112 27609 14176
rect 27673 14112 27689 14176
rect 27753 14112 27769 14176
rect 27833 14112 27849 14176
rect 27913 14112 27921 14176
rect 27601 13088 27921 14112
rect 27601 13024 27609 13088
rect 27673 13024 27689 13088
rect 27753 13024 27769 13088
rect 27833 13024 27849 13088
rect 27913 13024 27921 13088
rect 27601 12000 27921 13024
rect 27601 11936 27609 12000
rect 27673 11936 27689 12000
rect 27753 11936 27769 12000
rect 27833 11936 27849 12000
rect 27913 11936 27921 12000
rect 27601 10912 27921 11936
rect 27601 10848 27609 10912
rect 27673 10848 27689 10912
rect 27753 10848 27769 10912
rect 27833 10848 27849 10912
rect 27913 10848 27921 10912
rect 27601 9824 27921 10848
rect 27601 9760 27609 9824
rect 27673 9760 27689 9824
rect 27753 9760 27769 9824
rect 27833 9760 27849 9824
rect 27913 9760 27921 9824
rect 27601 8736 27921 9760
rect 27601 8672 27609 8736
rect 27673 8672 27689 8736
rect 27753 8672 27769 8736
rect 27833 8672 27849 8736
rect 27913 8672 27921 8736
rect 27601 7648 27921 8672
rect 27601 7584 27609 7648
rect 27673 7584 27689 7648
rect 27753 7584 27769 7648
rect 27833 7584 27849 7648
rect 27913 7584 27921 7648
rect 27601 6560 27921 7584
rect 27601 6496 27609 6560
rect 27673 6496 27689 6560
rect 27753 6496 27769 6560
rect 27833 6496 27849 6560
rect 27913 6496 27921 6560
rect 27601 5472 27921 6496
rect 27601 5408 27609 5472
rect 27673 5408 27689 5472
rect 27753 5408 27769 5472
rect 27833 5408 27849 5472
rect 27913 5408 27921 5472
rect 27601 4384 27921 5408
rect 27601 4320 27609 4384
rect 27673 4320 27689 4384
rect 27753 4320 27769 4384
rect 27833 4320 27849 4384
rect 27913 4320 27921 4384
rect 27601 3296 27921 4320
rect 27601 3232 27609 3296
rect 27673 3232 27689 3296
rect 27753 3232 27769 3296
rect 27833 3232 27849 3296
rect 27913 3232 27921 3296
rect 27601 2208 27921 3232
rect 27601 2144 27609 2208
rect 27673 2144 27689 2208
rect 27753 2144 27769 2208
rect 27833 2144 27849 2208
rect 27913 2144 27921 2208
rect 27601 1120 27921 2144
rect 27601 1056 27609 1120
rect 27673 1056 27689 1120
rect 27753 1056 27769 1120
rect 27833 1056 27849 1120
rect 27913 1056 27921 1120
rect 27601 496 27921 1056
rect 31488 21248 31808 21808
rect 31488 21184 31496 21248
rect 31560 21184 31576 21248
rect 31640 21184 31656 21248
rect 31720 21184 31736 21248
rect 31800 21184 31808 21248
rect 31488 20160 31808 21184
rect 31488 20096 31496 20160
rect 31560 20096 31576 20160
rect 31640 20096 31656 20160
rect 31720 20096 31736 20160
rect 31800 20096 31808 20160
rect 31488 19072 31808 20096
rect 31488 19008 31496 19072
rect 31560 19008 31576 19072
rect 31640 19008 31656 19072
rect 31720 19008 31736 19072
rect 31800 19008 31808 19072
rect 31488 17984 31808 19008
rect 31488 17920 31496 17984
rect 31560 17920 31576 17984
rect 31640 17920 31656 17984
rect 31720 17920 31736 17984
rect 31800 17920 31808 17984
rect 31488 16896 31808 17920
rect 31488 16832 31496 16896
rect 31560 16832 31576 16896
rect 31640 16832 31656 16896
rect 31720 16832 31736 16896
rect 31800 16832 31808 16896
rect 31488 15808 31808 16832
rect 31488 15744 31496 15808
rect 31560 15744 31576 15808
rect 31640 15744 31656 15808
rect 31720 15744 31736 15808
rect 31800 15744 31808 15808
rect 31488 14720 31808 15744
rect 31488 14656 31496 14720
rect 31560 14656 31576 14720
rect 31640 14656 31656 14720
rect 31720 14656 31736 14720
rect 31800 14656 31808 14720
rect 31488 13632 31808 14656
rect 31488 13568 31496 13632
rect 31560 13568 31576 13632
rect 31640 13568 31656 13632
rect 31720 13568 31736 13632
rect 31800 13568 31808 13632
rect 31488 12544 31808 13568
rect 31488 12480 31496 12544
rect 31560 12480 31576 12544
rect 31640 12480 31656 12544
rect 31720 12480 31736 12544
rect 31800 12480 31808 12544
rect 31488 11456 31808 12480
rect 31488 11392 31496 11456
rect 31560 11392 31576 11456
rect 31640 11392 31656 11456
rect 31720 11392 31736 11456
rect 31800 11392 31808 11456
rect 31488 10368 31808 11392
rect 31488 10304 31496 10368
rect 31560 10304 31576 10368
rect 31640 10304 31656 10368
rect 31720 10304 31736 10368
rect 31800 10304 31808 10368
rect 31488 9280 31808 10304
rect 31488 9216 31496 9280
rect 31560 9216 31576 9280
rect 31640 9216 31656 9280
rect 31720 9216 31736 9280
rect 31800 9216 31808 9280
rect 31488 8192 31808 9216
rect 31488 8128 31496 8192
rect 31560 8128 31576 8192
rect 31640 8128 31656 8192
rect 31720 8128 31736 8192
rect 31800 8128 31808 8192
rect 31488 7104 31808 8128
rect 31488 7040 31496 7104
rect 31560 7040 31576 7104
rect 31640 7040 31656 7104
rect 31720 7040 31736 7104
rect 31800 7040 31808 7104
rect 31488 6016 31808 7040
rect 31488 5952 31496 6016
rect 31560 5952 31576 6016
rect 31640 5952 31656 6016
rect 31720 5952 31736 6016
rect 31800 5952 31808 6016
rect 31488 4928 31808 5952
rect 31488 4864 31496 4928
rect 31560 4864 31576 4928
rect 31640 4864 31656 4928
rect 31720 4864 31736 4928
rect 31800 4864 31808 4928
rect 31488 3840 31808 4864
rect 31488 3776 31496 3840
rect 31560 3776 31576 3840
rect 31640 3776 31656 3840
rect 31720 3776 31736 3840
rect 31800 3776 31808 3840
rect 31488 2752 31808 3776
rect 31488 2688 31496 2752
rect 31560 2688 31576 2752
rect 31640 2688 31656 2752
rect 31720 2688 31736 2752
rect 31800 2688 31808 2752
rect 31488 1664 31808 2688
rect 31488 1600 31496 1664
rect 31560 1600 31576 1664
rect 31640 1600 31656 1664
rect 31720 1600 31736 1664
rect 31800 1600 31808 1664
rect 31488 576 31808 1600
rect 31488 512 31496 576
rect 31560 512 31576 576
rect 31640 512 31656 576
rect 31720 512 31736 576
rect 31800 512 31808 576
rect 31488 496 31808 512
use sky130_fd_sc_hd__and2_1  _01_
timestamp 0
transform -1 0 27232 0 1 21216
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _02_
timestamp 0
transform -1 0 26128 0 1 21216
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_3
timestamp 0
transform 1 0 828 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_15
timestamp 0
transform 1 0 1932 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_27
timestamp 0
transform 1 0 3036 0 1 544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_29
timestamp 0
transform 1 0 3220 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_41
timestamp 0
transform 1 0 4324 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_53
timestamp 0
transform 1 0 5428 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_57
timestamp 0
transform 1 0 5796 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_69
timestamp 0
transform 1 0 6900 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_81
timestamp 0
transform 1 0 8004 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_85
timestamp 0
transform 1 0 8372 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_97
timestamp 0
transform 1 0 9476 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_109
timestamp 0
transform 1 0 10580 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_113
timestamp 0
transform 1 0 10948 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_125
timestamp 0
transform 1 0 12052 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_137
timestamp 0
transform 1 0 13156 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_141
timestamp 0
transform 1 0 13524 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_153
timestamp 0
transform 1 0 14628 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_165
timestamp 0
transform 1 0 15732 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_169
timestamp 0
transform 1 0 16100 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_181
timestamp 0
transform 1 0 17204 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_193
timestamp 0
transform 1 0 18308 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_197
timestamp 0
transform 1 0 18676 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_209
timestamp 0
transform 1 0 19780 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_221
timestamp 0
transform 1 0 20884 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_225
timestamp 0
transform 1 0 21252 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_237
timestamp 0
transform 1 0 22356 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_249
timestamp 0
transform 1 0 23460 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_253
timestamp 0
transform 1 0 23828 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_265
timestamp 0
transform 1 0 24932 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_277
timestamp 0
transform 1 0 26036 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_281
timestamp 0
transform 1 0 26404 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_293
timestamp 0
transform 1 0 27508 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_305
timestamp 0
transform 1 0 28612 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_309
timestamp 0
transform 1 0 28980 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_321
timestamp 0
transform 1 0 30084 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_333
timestamp 0
transform 1 0 31188 0 1 544
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_3
timestamp 0
transform 1 0 828 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_15
timestamp 0
transform 1 0 1932 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_27
timestamp 0
transform 1 0 3036 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_39
timestamp 0
transform 1 0 4140 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_51
timestamp 0
transform 1 0 5244 0 -1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_55
timestamp 0
transform 1 0 5612 0 -1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_57
timestamp 0
transform 1 0 5796 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_69
timestamp 0
transform 1 0 6900 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_81
timestamp 0
transform 1 0 8004 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_93
timestamp 0
transform 1 0 9108 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_105
timestamp 0
transform 1 0 10212 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_111
timestamp 0
transform 1 0 10764 0 -1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_113
timestamp 0
transform 1 0 10948 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_125
timestamp 0
transform 1 0 12052 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_137
timestamp 0
transform 1 0 13156 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_149
timestamp 0
transform 1 0 14260 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_161
timestamp 0
transform 1 0 15364 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_167
timestamp 0
transform 1 0 15916 0 -1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_169
timestamp 0
transform 1 0 16100 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_181
timestamp 0
transform 1 0 17204 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_193
timestamp 0
transform 1 0 18308 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_205
timestamp 0
transform 1 0 19412 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_217
timestamp 0
transform 1 0 20516 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_223
timestamp 0
transform 1 0 21068 0 -1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_225
timestamp 0
transform 1 0 21252 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_237
timestamp 0
transform 1 0 22356 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_249
timestamp 0
transform 1 0 23460 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_261
timestamp 0
transform 1 0 24564 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_273
timestamp 0
transform 1 0 25668 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_279
timestamp 0
transform 1 0 26220 0 -1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_281
timestamp 0
transform 1 0 26404 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_293
timestamp 0
transform 1 0 27508 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_305
timestamp 0
transform 1 0 28612 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_317
timestamp 0
transform 1 0 29716 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_329
timestamp 0
transform 1 0 30820 0 -1 1632
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_3
timestamp 0
transform 1 0 828 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_15
timestamp 0
transform 1 0 1932 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 0
transform 1 0 3036 0 1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_29
timestamp 0
transform 1 0 3220 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_41
timestamp 0
transform 1 0 4324 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_53
timestamp 0
transform 1 0 5428 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_65
timestamp 0
transform 1 0 6532 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_77
timestamp 0
transform 1 0 7636 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_83
timestamp 0
transform 1 0 8188 0 1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_85
timestamp 0
transform 1 0 8372 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_97
timestamp 0
transform 1 0 9476 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_109
timestamp 0
transform 1 0 10580 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_121
timestamp 0
transform 1 0 11684 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_133
timestamp 0
transform 1 0 12788 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_139
timestamp 0
transform 1 0 13340 0 1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_141
timestamp 0
transform 1 0 13524 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_153
timestamp 0
transform 1 0 14628 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_165
timestamp 0
transform 1 0 15732 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_177
timestamp 0
transform 1 0 16836 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_189
timestamp 0
transform 1 0 17940 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_195
timestamp 0
transform 1 0 18492 0 1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_197
timestamp 0
transform 1 0 18676 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_209
timestamp 0
transform 1 0 19780 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_221
timestamp 0
transform 1 0 20884 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_233
timestamp 0
transform 1 0 21988 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_245
timestamp 0
transform 1 0 23092 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_251
timestamp 0
transform 1 0 23644 0 1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_253
timestamp 0
transform 1 0 23828 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_265
timestamp 0
transform 1 0 24932 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_277
timestamp 0
transform 1 0 26036 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_289
timestamp 0
transform 1 0 27140 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_301
timestamp 0
transform 1 0 28244 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_307
timestamp 0
transform 1 0 28796 0 1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_309
timestamp 0
transform 1 0 28980 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_321
timestamp 0
transform 1 0 30084 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_333
timestamp 0
transform 1 0 31188 0 1 1632
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_3
timestamp 0
transform 1 0 828 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_15
timestamp 0
transform 1 0 1932 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_27
timestamp 0
transform 1 0 3036 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_39
timestamp 0
transform 1 0 4140 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_51
timestamp 0
transform 1 0 5244 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_55
timestamp 0
transform 1 0 5612 0 -1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_57
timestamp 0
transform 1 0 5796 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_69
timestamp 0
transform 1 0 6900 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_81
timestamp 0
transform 1 0 8004 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_93
timestamp 0
transform 1 0 9108 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_105
timestamp 0
transform 1 0 10212 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_111
timestamp 0
transform 1 0 10764 0 -1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_113
timestamp 0
transform 1 0 10948 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_125
timestamp 0
transform 1 0 12052 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_137
timestamp 0
transform 1 0 13156 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_149
timestamp 0
transform 1 0 14260 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_161
timestamp 0
transform 1 0 15364 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_167
timestamp 0
transform 1 0 15916 0 -1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_169
timestamp 0
transform 1 0 16100 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_181
timestamp 0
transform 1 0 17204 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_193
timestamp 0
transform 1 0 18308 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_205
timestamp 0
transform 1 0 19412 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_217
timestamp 0
transform 1 0 20516 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_223
timestamp 0
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_225
timestamp 0
transform 1 0 21252 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_237
timestamp 0
transform 1 0 22356 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_249
timestamp 0
transform 1 0 23460 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_261
timestamp 0
transform 1 0 24564 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_273
timestamp 0
transform 1 0 25668 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_279
timestamp 0
transform 1 0 26220 0 -1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_281
timestamp 0
transform 1 0 26404 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_293
timestamp 0
transform 1 0 27508 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_305
timestamp 0
transform 1 0 28612 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_317
timestamp 0
transform 1 0 29716 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_329
timestamp 0
transform 1 0 30820 0 -1 2720
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_3
timestamp 0
transform 1 0 828 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_15
timestamp 0
transform 1 0 1932 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp 0
transform 1 0 3036 0 1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_29
timestamp 0
transform 1 0 3220 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_41
timestamp 0
transform 1 0 4324 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_53
timestamp 0
transform 1 0 5428 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_65
timestamp 0
transform 1 0 6532 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_77
timestamp 0
transform 1 0 7636 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_83
timestamp 0
transform 1 0 8188 0 1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_85
timestamp 0
transform 1 0 8372 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_97
timestamp 0
transform 1 0 9476 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_109
timestamp 0
transform 1 0 10580 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_121
timestamp 0
transform 1 0 11684 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_133
timestamp 0
transform 1 0 12788 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_139
timestamp 0
transform 1 0 13340 0 1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_141
timestamp 0
transform 1 0 13524 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_153
timestamp 0
transform 1 0 14628 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_165
timestamp 0
transform 1 0 15732 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_177
timestamp 0
transform 1 0 16836 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_189
timestamp 0
transform 1 0 17940 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_195
timestamp 0
transform 1 0 18492 0 1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_197
timestamp 0
transform 1 0 18676 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_209
timestamp 0
transform 1 0 19780 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_221
timestamp 0
transform 1 0 20884 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_233
timestamp 0
transform 1 0 21988 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_245
timestamp 0
transform 1 0 23092 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_251
timestamp 0
transform 1 0 23644 0 1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_253
timestamp 0
transform 1 0 23828 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_265
timestamp 0
transform 1 0 24932 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_277
timestamp 0
transform 1 0 26036 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_289
timestamp 0
transform 1 0 27140 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_301
timestamp 0
transform 1 0 28244 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_307
timestamp 0
transform 1 0 28796 0 1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_309
timestamp 0
transform 1 0 28980 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_321
timestamp 0
transform 1 0 30084 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_333
timestamp 0
transform 1 0 31188 0 1 2720
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_3
timestamp 0
transform 1 0 828 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_15
timestamp 0
transform 1 0 1932 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_27
timestamp 0
transform 1 0 3036 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_39
timestamp 0
transform 1 0 4140 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_51
timestamp 0
transform 1 0 5244 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_55
timestamp 0
transform 1 0 5612 0 -1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_57
timestamp 0
transform 1 0 5796 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_69
timestamp 0
transform 1 0 6900 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_81
timestamp 0
transform 1 0 8004 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_93
timestamp 0
transform 1 0 9108 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_105
timestamp 0
transform 1 0 10212 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_111
timestamp 0
transform 1 0 10764 0 -1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_113
timestamp 0
transform 1 0 10948 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_125
timestamp 0
transform 1 0 12052 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_137
timestamp 0
transform 1 0 13156 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_149
timestamp 0
transform 1 0 14260 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_161
timestamp 0
transform 1 0 15364 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_167
timestamp 0
transform 1 0 15916 0 -1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_169
timestamp 0
transform 1 0 16100 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_181
timestamp 0
transform 1 0 17204 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_193
timestamp 0
transform 1 0 18308 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_205
timestamp 0
transform 1 0 19412 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_217
timestamp 0
transform 1 0 20516 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_223
timestamp 0
transform 1 0 21068 0 -1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_225
timestamp 0
transform 1 0 21252 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_237
timestamp 0
transform 1 0 22356 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_249
timestamp 0
transform 1 0 23460 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_261
timestamp 0
transform 1 0 24564 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_273
timestamp 0
transform 1 0 25668 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_279
timestamp 0
transform 1 0 26220 0 -1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_281
timestamp 0
transform 1 0 26404 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_293
timestamp 0
transform 1 0 27508 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_305
timestamp 0
transform 1 0 28612 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_317
timestamp 0
transform 1 0 29716 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_329
timestamp 0
transform 1 0 30820 0 -1 3808
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_3
timestamp 0
transform 1 0 828 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_15
timestamp 0
transform 1 0 1932 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_27
timestamp 0
transform 1 0 3036 0 1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_29
timestamp 0
transform 1 0 3220 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_41
timestamp 0
transform 1 0 4324 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_53
timestamp 0
transform 1 0 5428 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_65
timestamp 0
transform 1 0 6532 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_77
timestamp 0
transform 1 0 7636 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_83
timestamp 0
transform 1 0 8188 0 1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_85
timestamp 0
transform 1 0 8372 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_97
timestamp 0
transform 1 0 9476 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_109
timestamp 0
transform 1 0 10580 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_121
timestamp 0
transform 1 0 11684 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_133
timestamp 0
transform 1 0 12788 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_139
timestamp 0
transform 1 0 13340 0 1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_141
timestamp 0
transform 1 0 13524 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_153
timestamp 0
transform 1 0 14628 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_165
timestamp 0
transform 1 0 15732 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_177
timestamp 0
transform 1 0 16836 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_189
timestamp 0
transform 1 0 17940 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_195
timestamp 0
transform 1 0 18492 0 1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_197
timestamp 0
transform 1 0 18676 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_209
timestamp 0
transform 1 0 19780 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_221
timestamp 0
transform 1 0 20884 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_233
timestamp 0
transform 1 0 21988 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_245
timestamp 0
transform 1 0 23092 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_251
timestamp 0
transform 1 0 23644 0 1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_253
timestamp 0
transform 1 0 23828 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_265
timestamp 0
transform 1 0 24932 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_277
timestamp 0
transform 1 0 26036 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_289
timestamp 0
transform 1 0 27140 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_301
timestamp 0
transform 1 0 28244 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_307
timestamp 0
transform 1 0 28796 0 1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_309
timestamp 0
transform 1 0 28980 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_321
timestamp 0
transform 1 0 30084 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_333
timestamp 0
transform 1 0 31188 0 1 3808
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_3
timestamp 0
transform 1 0 828 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_15
timestamp 0
transform 1 0 1932 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_27
timestamp 0
transform 1 0 3036 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_39
timestamp 0
transform 1 0 4140 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_51
timestamp 0
transform 1 0 5244 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_55
timestamp 0
transform 1 0 5612 0 -1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_57
timestamp 0
transform 1 0 5796 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_69
timestamp 0
transform 1 0 6900 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_81
timestamp 0
transform 1 0 8004 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_93
timestamp 0
transform 1 0 9108 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_105
timestamp 0
transform 1 0 10212 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_111
timestamp 0
transform 1 0 10764 0 -1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_113
timestamp 0
transform 1 0 10948 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_125
timestamp 0
transform 1 0 12052 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_137
timestamp 0
transform 1 0 13156 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_149
timestamp 0
transform 1 0 14260 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_161
timestamp 0
transform 1 0 15364 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_167
timestamp 0
transform 1 0 15916 0 -1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_169
timestamp 0
transform 1 0 16100 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_181
timestamp 0
transform 1 0 17204 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_193
timestamp 0
transform 1 0 18308 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_205
timestamp 0
transform 1 0 19412 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_217
timestamp 0
transform 1 0 20516 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_223
timestamp 0
transform 1 0 21068 0 -1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_225
timestamp 0
transform 1 0 21252 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_237
timestamp 0
transform 1 0 22356 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_249
timestamp 0
transform 1 0 23460 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_261
timestamp 0
transform 1 0 24564 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_273
timestamp 0
transform 1 0 25668 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_279
timestamp 0
transform 1 0 26220 0 -1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_281
timestamp 0
transform 1 0 26404 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_293
timestamp 0
transform 1 0 27508 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_305
timestamp 0
transform 1 0 28612 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_317
timestamp 0
transform 1 0 29716 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_329
timestamp 0
transform 1 0 30820 0 -1 4896
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_3
timestamp 0
transform 1 0 828 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_15
timestamp 0
transform 1 0 1932 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_27
timestamp 0
transform 1 0 3036 0 1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_29
timestamp 0
transform 1 0 3220 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_41
timestamp 0
transform 1 0 4324 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_53
timestamp 0
transform 1 0 5428 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_65
timestamp 0
transform 1 0 6532 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_77
timestamp 0
transform 1 0 7636 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_83
timestamp 0
transform 1 0 8188 0 1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_85
timestamp 0
transform 1 0 8372 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_97
timestamp 0
transform 1 0 9476 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_109
timestamp 0
transform 1 0 10580 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_121
timestamp 0
transform 1 0 11684 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_133
timestamp 0
transform 1 0 12788 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_139
timestamp 0
transform 1 0 13340 0 1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_141
timestamp 0
transform 1 0 13524 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_153
timestamp 0
transform 1 0 14628 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_165
timestamp 0
transform 1 0 15732 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_177
timestamp 0
transform 1 0 16836 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_189
timestamp 0
transform 1 0 17940 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_195
timestamp 0
transform 1 0 18492 0 1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_197
timestamp 0
transform 1 0 18676 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_209
timestamp 0
transform 1 0 19780 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_221
timestamp 0
transform 1 0 20884 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_233
timestamp 0
transform 1 0 21988 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_245
timestamp 0
transform 1 0 23092 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_251
timestamp 0
transform 1 0 23644 0 1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_253
timestamp 0
transform 1 0 23828 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_265
timestamp 0
transform 1 0 24932 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_277
timestamp 0
transform 1 0 26036 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_289
timestamp 0
transform 1 0 27140 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_301
timestamp 0
transform 1 0 28244 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_307
timestamp 0
transform 1 0 28796 0 1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_309
timestamp 0
transform 1 0 28980 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_321
timestamp 0
transform 1 0 30084 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_333
timestamp 0
transform 1 0 31188 0 1 4896
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_3
timestamp 0
transform 1 0 828 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_15
timestamp 0
transform 1 0 1932 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_27
timestamp 0
transform 1 0 3036 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_39
timestamp 0
transform 1 0 4140 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_51
timestamp 0
transform 1 0 5244 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_55
timestamp 0
transform 1 0 5612 0 -1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_57
timestamp 0
transform 1 0 5796 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_69
timestamp 0
transform 1 0 6900 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_81
timestamp 0
transform 1 0 8004 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_93
timestamp 0
transform 1 0 9108 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_105
timestamp 0
transform 1 0 10212 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_111
timestamp 0
transform 1 0 10764 0 -1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_113
timestamp 0
transform 1 0 10948 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_125
timestamp 0
transform 1 0 12052 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_137
timestamp 0
transform 1 0 13156 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_149
timestamp 0
transform 1 0 14260 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_161
timestamp 0
transform 1 0 15364 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_167
timestamp 0
transform 1 0 15916 0 -1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_169
timestamp 0
transform 1 0 16100 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_181
timestamp 0
transform 1 0 17204 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_193
timestamp 0
transform 1 0 18308 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_205
timestamp 0
transform 1 0 19412 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_217
timestamp 0
transform 1 0 20516 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_223
timestamp 0
transform 1 0 21068 0 -1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_225
timestamp 0
transform 1 0 21252 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_237
timestamp 0
transform 1 0 22356 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_249
timestamp 0
transform 1 0 23460 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_261
timestamp 0
transform 1 0 24564 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_273
timestamp 0
transform 1 0 25668 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_279
timestamp 0
transform 1 0 26220 0 -1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_281
timestamp 0
transform 1 0 26404 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_293
timestamp 0
transform 1 0 27508 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_305
timestamp 0
transform 1 0 28612 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_317
timestamp 0
transform 1 0 29716 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_329
timestamp 0
transform 1 0 30820 0 -1 5984
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_3
timestamp 0
transform 1 0 828 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_15
timestamp 0
transform 1 0 1932 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_27
timestamp 0
transform 1 0 3036 0 1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_29
timestamp 0
transform 1 0 3220 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_41
timestamp 0
transform 1 0 4324 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_53
timestamp 0
transform 1 0 5428 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_65
timestamp 0
transform 1 0 6532 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_77
timestamp 0
transform 1 0 7636 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_83
timestamp 0
transform 1 0 8188 0 1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_85
timestamp 0
transform 1 0 8372 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_97
timestamp 0
transform 1 0 9476 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_109
timestamp 0
transform 1 0 10580 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_121
timestamp 0
transform 1 0 11684 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_133
timestamp 0
transform 1 0 12788 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_139
timestamp 0
transform 1 0 13340 0 1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_141
timestamp 0
transform 1 0 13524 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_153
timestamp 0
transform 1 0 14628 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_165
timestamp 0
transform 1 0 15732 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_177
timestamp 0
transform 1 0 16836 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_189
timestamp 0
transform 1 0 17940 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_195
timestamp 0
transform 1 0 18492 0 1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_197
timestamp 0
transform 1 0 18676 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_209
timestamp 0
transform 1 0 19780 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_221
timestamp 0
transform 1 0 20884 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_233
timestamp 0
transform 1 0 21988 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_245
timestamp 0
transform 1 0 23092 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_251
timestamp 0
transform 1 0 23644 0 1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_253
timestamp 0
transform 1 0 23828 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_265
timestamp 0
transform 1 0 24932 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_277
timestamp 0
transform 1 0 26036 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_289
timestamp 0
transform 1 0 27140 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_301
timestamp 0
transform 1 0 28244 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_307
timestamp 0
transform 1 0 28796 0 1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_309
timestamp 0
transform 1 0 28980 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_321
timestamp 0
transform 1 0 30084 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_333
timestamp 0
transform 1 0 31188 0 1 5984
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_3
timestamp 0
transform 1 0 828 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_15
timestamp 0
transform 1 0 1932 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_27
timestamp 0
transform 1 0 3036 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_39
timestamp 0
transform 1 0 4140 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_51
timestamp 0
transform 1 0 5244 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_55
timestamp 0
transform 1 0 5612 0 -1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_57
timestamp 0
transform 1 0 5796 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_69
timestamp 0
transform 1 0 6900 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_81
timestamp 0
transform 1 0 8004 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_93
timestamp 0
transform 1 0 9108 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_105
timestamp 0
transform 1 0 10212 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_111
timestamp 0
transform 1 0 10764 0 -1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_113
timestamp 0
transform 1 0 10948 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_125
timestamp 0
transform 1 0 12052 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_137
timestamp 0
transform 1 0 13156 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_149
timestamp 0
transform 1 0 14260 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_161
timestamp 0
transform 1 0 15364 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_167
timestamp 0
transform 1 0 15916 0 -1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_169
timestamp 0
transform 1 0 16100 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_181
timestamp 0
transform 1 0 17204 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_193
timestamp 0
transform 1 0 18308 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_205
timestamp 0
transform 1 0 19412 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_217
timestamp 0
transform 1 0 20516 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_223
timestamp 0
transform 1 0 21068 0 -1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_225
timestamp 0
transform 1 0 21252 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_237
timestamp 0
transform 1 0 22356 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_249
timestamp 0
transform 1 0 23460 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_261
timestamp 0
transform 1 0 24564 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_273
timestamp 0
transform 1 0 25668 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_279
timestamp 0
transform 1 0 26220 0 -1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_281
timestamp 0
transform 1 0 26404 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_293
timestamp 0
transform 1 0 27508 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_305
timestamp 0
transform 1 0 28612 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_317
timestamp 0
transform 1 0 29716 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_329
timestamp 0
transform 1 0 30820 0 -1 7072
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_3
timestamp 0
transform 1 0 828 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_15
timestamp 0
transform 1 0 1932 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_27
timestamp 0
transform 1 0 3036 0 1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_29
timestamp 0
transform 1 0 3220 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_41
timestamp 0
transform 1 0 4324 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_53
timestamp 0
transform 1 0 5428 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_65
timestamp 0
transform 1 0 6532 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_77
timestamp 0
transform 1 0 7636 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_83
timestamp 0
transform 1 0 8188 0 1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_85
timestamp 0
transform 1 0 8372 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_97
timestamp 0
transform 1 0 9476 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_109
timestamp 0
transform 1 0 10580 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_121
timestamp 0
transform 1 0 11684 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_133
timestamp 0
transform 1 0 12788 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_139
timestamp 0
transform 1 0 13340 0 1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_141
timestamp 0
transform 1 0 13524 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_153
timestamp 0
transform 1 0 14628 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_165
timestamp 0
transform 1 0 15732 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_177
timestamp 0
transform 1 0 16836 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_189
timestamp 0
transform 1 0 17940 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_195
timestamp 0
transform 1 0 18492 0 1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_197
timestamp 0
transform 1 0 18676 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_209
timestamp 0
transform 1 0 19780 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_221
timestamp 0
transform 1 0 20884 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_233
timestamp 0
transform 1 0 21988 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_245
timestamp 0
transform 1 0 23092 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_251
timestamp 0
transform 1 0 23644 0 1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_253
timestamp 0
transform 1 0 23828 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_265
timestamp 0
transform 1 0 24932 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_277
timestamp 0
transform 1 0 26036 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_289
timestamp 0
transform 1 0 27140 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_301
timestamp 0
transform 1 0 28244 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_307
timestamp 0
transform 1 0 28796 0 1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_309
timestamp 0
transform 1 0 28980 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_321
timestamp 0
transform 1 0 30084 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_333
timestamp 0
transform 1 0 31188 0 1 7072
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_3
timestamp 0
transform 1 0 828 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_15
timestamp 0
transform 1 0 1932 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_27
timestamp 0
transform 1 0 3036 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_39
timestamp 0
transform 1 0 4140 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_51
timestamp 0
transform 1 0 5244 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_55
timestamp 0
transform 1 0 5612 0 -1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_57
timestamp 0
transform 1 0 5796 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_69
timestamp 0
transform 1 0 6900 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_81
timestamp 0
transform 1 0 8004 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_93
timestamp 0
transform 1 0 9108 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_105
timestamp 0
transform 1 0 10212 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_111
timestamp 0
transform 1 0 10764 0 -1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_113
timestamp 0
transform 1 0 10948 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_125
timestamp 0
transform 1 0 12052 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_137
timestamp 0
transform 1 0 13156 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_149
timestamp 0
transform 1 0 14260 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_161
timestamp 0
transform 1 0 15364 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_167
timestamp 0
transform 1 0 15916 0 -1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_169
timestamp 0
transform 1 0 16100 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_181
timestamp 0
transform 1 0 17204 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_193
timestamp 0
transform 1 0 18308 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_205
timestamp 0
transform 1 0 19412 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_217
timestamp 0
transform 1 0 20516 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_223
timestamp 0
transform 1 0 21068 0 -1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_225
timestamp 0
transform 1 0 21252 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_237
timestamp 0
transform 1 0 22356 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_249
timestamp 0
transform 1 0 23460 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_261
timestamp 0
transform 1 0 24564 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_273
timestamp 0
transform 1 0 25668 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_279
timestamp 0
transform 1 0 26220 0 -1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_281
timestamp 0
transform 1 0 26404 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_293
timestamp 0
transform 1 0 27508 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_305
timestamp 0
transform 1 0 28612 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_317
timestamp 0
transform 1 0 29716 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_329
timestamp 0
transform 1 0 30820 0 -1 8160
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_3
timestamp 0
transform 1 0 828 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_15
timestamp 0
transform 1 0 1932 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_27
timestamp 0
transform 1 0 3036 0 1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_29
timestamp 0
transform 1 0 3220 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_41
timestamp 0
transform 1 0 4324 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_53
timestamp 0
transform 1 0 5428 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_65
timestamp 0
transform 1 0 6532 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_77
timestamp 0
transform 1 0 7636 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_83
timestamp 0
transform 1 0 8188 0 1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_85
timestamp 0
transform 1 0 8372 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_97
timestamp 0
transform 1 0 9476 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_109
timestamp 0
transform 1 0 10580 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_121
timestamp 0
transform 1 0 11684 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_133
timestamp 0
transform 1 0 12788 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_139
timestamp 0
transform 1 0 13340 0 1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_141
timestamp 0
transform 1 0 13524 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_153
timestamp 0
transform 1 0 14628 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_165
timestamp 0
transform 1 0 15732 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_177
timestamp 0
transform 1 0 16836 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_189
timestamp 0
transform 1 0 17940 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_195
timestamp 0
transform 1 0 18492 0 1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_197
timestamp 0
transform 1 0 18676 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_209
timestamp 0
transform 1 0 19780 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_221
timestamp 0
transform 1 0 20884 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_233
timestamp 0
transform 1 0 21988 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_245
timestamp 0
transform 1 0 23092 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_251
timestamp 0
transform 1 0 23644 0 1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_253
timestamp 0
transform 1 0 23828 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_265
timestamp 0
transform 1 0 24932 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_277
timestamp 0
transform 1 0 26036 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_289
timestamp 0
transform 1 0 27140 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_301
timestamp 0
transform 1 0 28244 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_307
timestamp 0
transform 1 0 28796 0 1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_309
timestamp 0
transform 1 0 28980 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_321
timestamp 0
transform 1 0 30084 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_333
timestamp 0
transform 1 0 31188 0 1 8160
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_3
timestamp 0
transform 1 0 828 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_15
timestamp 0
transform 1 0 1932 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_27
timestamp 0
transform 1 0 3036 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_39
timestamp 0
transform 1 0 4140 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_51
timestamp 0
transform 1 0 5244 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_55
timestamp 0
transform 1 0 5612 0 -1 9248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_57
timestamp 0
transform 1 0 5796 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_69
timestamp 0
transform 1 0 6900 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_81
timestamp 0
transform 1 0 8004 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_93
timestamp 0
transform 1 0 9108 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_105
timestamp 0
transform 1 0 10212 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_111
timestamp 0
transform 1 0 10764 0 -1 9248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_113
timestamp 0
transform 1 0 10948 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_125
timestamp 0
transform 1 0 12052 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_137
timestamp 0
transform 1 0 13156 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_149
timestamp 0
transform 1 0 14260 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_161
timestamp 0
transform 1 0 15364 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_167
timestamp 0
transform 1 0 15916 0 -1 9248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_169
timestamp 0
transform 1 0 16100 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_181
timestamp 0
transform 1 0 17204 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_193
timestamp 0
transform 1 0 18308 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_205
timestamp 0
transform 1 0 19412 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_217
timestamp 0
transform 1 0 20516 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_223
timestamp 0
transform 1 0 21068 0 -1 9248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_225
timestamp 0
transform 1 0 21252 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_237
timestamp 0
transform 1 0 22356 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_249
timestamp 0
transform 1 0 23460 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_261
timestamp 0
transform 1 0 24564 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_273
timestamp 0
transform 1 0 25668 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_279
timestamp 0
transform 1 0 26220 0 -1 9248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_281
timestamp 0
transform 1 0 26404 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_293
timestamp 0
transform 1 0 27508 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_305
timestamp 0
transform 1 0 28612 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_317
timestamp 0
transform 1 0 29716 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_329
timestamp 0
transform 1 0 30820 0 -1 9248
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_3
timestamp 0
transform 1 0 828 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_15
timestamp 0
transform 1 0 1932 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_27
timestamp 0
transform 1 0 3036 0 1 9248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_29
timestamp 0
transform 1 0 3220 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_41
timestamp 0
transform 1 0 4324 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_53
timestamp 0
transform 1 0 5428 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_65
timestamp 0
transform 1 0 6532 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_77
timestamp 0
transform 1 0 7636 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_83
timestamp 0
transform 1 0 8188 0 1 9248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_85
timestamp 0
transform 1 0 8372 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_97
timestamp 0
transform 1 0 9476 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_109
timestamp 0
transform 1 0 10580 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_121
timestamp 0
transform 1 0 11684 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_133
timestamp 0
transform 1 0 12788 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_139
timestamp 0
transform 1 0 13340 0 1 9248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_141
timestamp 0
transform 1 0 13524 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_153
timestamp 0
transform 1 0 14628 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_165
timestamp 0
transform 1 0 15732 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_177
timestamp 0
transform 1 0 16836 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_189
timestamp 0
transform 1 0 17940 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_195
timestamp 0
transform 1 0 18492 0 1 9248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_197
timestamp 0
transform 1 0 18676 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_209
timestamp 0
transform 1 0 19780 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_221
timestamp 0
transform 1 0 20884 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_233
timestamp 0
transform 1 0 21988 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_245
timestamp 0
transform 1 0 23092 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_251
timestamp 0
transform 1 0 23644 0 1 9248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_253
timestamp 0
transform 1 0 23828 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_265
timestamp 0
transform 1 0 24932 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_277
timestamp 0
transform 1 0 26036 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_289
timestamp 0
transform 1 0 27140 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_301
timestamp 0
transform 1 0 28244 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_307
timestamp 0
transform 1 0 28796 0 1 9248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_309
timestamp 0
transform 1 0 28980 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_321
timestamp 0
transform 1 0 30084 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_333
timestamp 0
transform 1 0 31188 0 1 9248
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_3
timestamp 0
transform 1 0 828 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_15
timestamp 0
transform 1 0 1932 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_27
timestamp 0
transform 1 0 3036 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_39
timestamp 0
transform 1 0 4140 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_51
timestamp 0
transform 1 0 5244 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_55
timestamp 0
transform 1 0 5612 0 -1 10336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_57
timestamp 0
transform 1 0 5796 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_69
timestamp 0
transform 1 0 6900 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_81
timestamp 0
transform 1 0 8004 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_93
timestamp 0
transform 1 0 9108 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_105
timestamp 0
transform 1 0 10212 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_111
timestamp 0
transform 1 0 10764 0 -1 10336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_113
timestamp 0
transform 1 0 10948 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_125
timestamp 0
transform 1 0 12052 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_137
timestamp 0
transform 1 0 13156 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_149
timestamp 0
transform 1 0 14260 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_161
timestamp 0
transform 1 0 15364 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_167
timestamp 0
transform 1 0 15916 0 -1 10336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_169
timestamp 0
transform 1 0 16100 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_181
timestamp 0
transform 1 0 17204 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_193
timestamp 0
transform 1 0 18308 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_205
timestamp 0
transform 1 0 19412 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_217
timestamp 0
transform 1 0 20516 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_223
timestamp 0
transform 1 0 21068 0 -1 10336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_225
timestamp 0
transform 1 0 21252 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_237
timestamp 0
transform 1 0 22356 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_249
timestamp 0
transform 1 0 23460 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_261
timestamp 0
transform 1 0 24564 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_273
timestamp 0
transform 1 0 25668 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_279
timestamp 0
transform 1 0 26220 0 -1 10336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_281
timestamp 0
transform 1 0 26404 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_293
timestamp 0
transform 1 0 27508 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_305
timestamp 0
transform 1 0 28612 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_317
timestamp 0
transform 1 0 29716 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_329
timestamp 0
transform 1 0 30820 0 -1 10336
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_3
timestamp 0
transform 1 0 828 0 1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_15
timestamp 0
transform 1 0 1932 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_27
timestamp 0
transform 1 0 3036 0 1 10336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_29
timestamp 0
transform 1 0 3220 0 1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_41
timestamp 0
transform 1 0 4324 0 1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_53
timestamp 0
transform 1 0 5428 0 1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_65
timestamp 0
transform 1 0 6532 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_77
timestamp 0
transform 1 0 7636 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_83
timestamp 0
transform 1 0 8188 0 1 10336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_85
timestamp 0
transform 1 0 8372 0 1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_97
timestamp 0
transform 1 0 9476 0 1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_109
timestamp 0
transform 1 0 10580 0 1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_121
timestamp 0
transform 1 0 11684 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_133
timestamp 0
transform 1 0 12788 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_139
timestamp 0
transform 1 0 13340 0 1 10336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_141
timestamp 0
transform 1 0 13524 0 1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_153
timestamp 0
transform 1 0 14628 0 1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_165
timestamp 0
transform 1 0 15732 0 1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_177
timestamp 0
transform 1 0 16836 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_189
timestamp 0
transform 1 0 17940 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_195
timestamp 0
transform 1 0 18492 0 1 10336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_197
timestamp 0
transform 1 0 18676 0 1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_209
timestamp 0
transform 1 0 19780 0 1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_221
timestamp 0
transform 1 0 20884 0 1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_233
timestamp 0
transform 1 0 21988 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_245
timestamp 0
transform 1 0 23092 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_251
timestamp 0
transform 1 0 23644 0 1 10336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_253
timestamp 0
transform 1 0 23828 0 1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_265
timestamp 0
transform 1 0 24932 0 1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_277
timestamp 0
transform 1 0 26036 0 1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_289
timestamp 0
transform 1 0 27140 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_301
timestamp 0
transform 1 0 28244 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_307
timestamp 0
transform 1 0 28796 0 1 10336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_309
timestamp 0
transform 1 0 28980 0 1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_321
timestamp 0
transform 1 0 30084 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_333
timestamp 0
transform 1 0 31188 0 1 10336
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_3
timestamp 0
transform 1 0 828 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_15
timestamp 0
transform 1 0 1932 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_27
timestamp 0
transform 1 0 3036 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_39
timestamp 0
transform 1 0 4140 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_51
timestamp 0
transform 1 0 5244 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_55
timestamp 0
transform 1 0 5612 0 -1 11424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_57
timestamp 0
transform 1 0 5796 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_69
timestamp 0
transform 1 0 6900 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_81
timestamp 0
transform 1 0 8004 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_93
timestamp 0
transform 1 0 9108 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_105
timestamp 0
transform 1 0 10212 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_111
timestamp 0
transform 1 0 10764 0 -1 11424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_113
timestamp 0
transform 1 0 10948 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_125
timestamp 0
transform 1 0 12052 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_137
timestamp 0
transform 1 0 13156 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_149
timestamp 0
transform 1 0 14260 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_161
timestamp 0
transform 1 0 15364 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_167
timestamp 0
transform 1 0 15916 0 -1 11424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_169
timestamp 0
transform 1 0 16100 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_181
timestamp 0
transform 1 0 17204 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_193
timestamp 0
transform 1 0 18308 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_205
timestamp 0
transform 1 0 19412 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_217
timestamp 0
transform 1 0 20516 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_223
timestamp 0
transform 1 0 21068 0 -1 11424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_225
timestamp 0
transform 1 0 21252 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_237
timestamp 0
transform 1 0 22356 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_249
timestamp 0
transform 1 0 23460 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_261
timestamp 0
transform 1 0 24564 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_273
timestamp 0
transform 1 0 25668 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_279
timestamp 0
transform 1 0 26220 0 -1 11424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_281
timestamp 0
transform 1 0 26404 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_293
timestamp 0
transform 1 0 27508 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_305
timestamp 0
transform 1 0 28612 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_317
timestamp 0
transform 1 0 29716 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_329
timestamp 0
transform 1 0 30820 0 -1 11424
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_3
timestamp 0
transform 1 0 828 0 1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_15
timestamp 0
transform 1 0 1932 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_27
timestamp 0
transform 1 0 3036 0 1 11424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_29
timestamp 0
transform 1 0 3220 0 1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_41
timestamp 0
transform 1 0 4324 0 1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_53
timestamp 0
transform 1 0 5428 0 1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_65
timestamp 0
transform 1 0 6532 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_77
timestamp 0
transform 1 0 7636 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_83
timestamp 0
transform 1 0 8188 0 1 11424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_85
timestamp 0
transform 1 0 8372 0 1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_97
timestamp 0
transform 1 0 9476 0 1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_109
timestamp 0
transform 1 0 10580 0 1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_121
timestamp 0
transform 1 0 11684 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_133
timestamp 0
transform 1 0 12788 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_139
timestamp 0
transform 1 0 13340 0 1 11424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_141
timestamp 0
transform 1 0 13524 0 1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_153
timestamp 0
transform 1 0 14628 0 1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_165
timestamp 0
transform 1 0 15732 0 1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_177
timestamp 0
transform 1 0 16836 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_189
timestamp 0
transform 1 0 17940 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_195
timestamp 0
transform 1 0 18492 0 1 11424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_197
timestamp 0
transform 1 0 18676 0 1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_209
timestamp 0
transform 1 0 19780 0 1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_221
timestamp 0
transform 1 0 20884 0 1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_233
timestamp 0
transform 1 0 21988 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_245
timestamp 0
transform 1 0 23092 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_251
timestamp 0
transform 1 0 23644 0 1 11424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_253
timestamp 0
transform 1 0 23828 0 1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_265
timestamp 0
transform 1 0 24932 0 1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_277
timestamp 0
transform 1 0 26036 0 1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_289
timestamp 0
transform 1 0 27140 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_301
timestamp 0
transform 1 0 28244 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_307
timestamp 0
transform 1 0 28796 0 1 11424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_309
timestamp 0
transform 1 0 28980 0 1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_321
timestamp 0
transform 1 0 30084 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_333
timestamp 0
transform 1 0 31188 0 1 11424
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_3
timestamp 0
transform 1 0 828 0 -1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_15
timestamp 0
transform 1 0 1932 0 -1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_27
timestamp 0
transform 1 0 3036 0 -1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_39
timestamp 0
transform 1 0 4140 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_51
timestamp 0
transform 1 0 5244 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_55
timestamp 0
transform 1 0 5612 0 -1 12512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_57
timestamp 0
transform 1 0 5796 0 -1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_69
timestamp 0
transform 1 0 6900 0 -1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_81
timestamp 0
transform 1 0 8004 0 -1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_93
timestamp 0
transform 1 0 9108 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_105
timestamp 0
transform 1 0 10212 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_111
timestamp 0
transform 1 0 10764 0 -1 12512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_113
timestamp 0
transform 1 0 10948 0 -1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_125
timestamp 0
transform 1 0 12052 0 -1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_137
timestamp 0
transform 1 0 13156 0 -1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_149
timestamp 0
transform 1 0 14260 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_161
timestamp 0
transform 1 0 15364 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_167
timestamp 0
transform 1 0 15916 0 -1 12512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_169
timestamp 0
transform 1 0 16100 0 -1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_181
timestamp 0
transform 1 0 17204 0 -1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_193
timestamp 0
transform 1 0 18308 0 -1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_205
timestamp 0
transform 1 0 19412 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_217
timestamp 0
transform 1 0 20516 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_223
timestamp 0
transform 1 0 21068 0 -1 12512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_225
timestamp 0
transform 1 0 21252 0 -1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_237
timestamp 0
transform 1 0 22356 0 -1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_249
timestamp 0
transform 1 0 23460 0 -1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_261
timestamp 0
transform 1 0 24564 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_273
timestamp 0
transform 1 0 25668 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_279
timestamp 0
transform 1 0 26220 0 -1 12512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_281
timestamp 0
transform 1 0 26404 0 -1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_293
timestamp 0
transform 1 0 27508 0 -1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_305
timestamp 0
transform 1 0 28612 0 -1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_317
timestamp 0
transform 1 0 29716 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_329
timestamp 0
transform 1 0 30820 0 -1 12512
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_3
timestamp 0
transform 1 0 828 0 1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_15
timestamp 0
transform 1 0 1932 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_27
timestamp 0
transform 1 0 3036 0 1 12512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_29
timestamp 0
transform 1 0 3220 0 1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_41
timestamp 0
transform 1 0 4324 0 1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_53
timestamp 0
transform 1 0 5428 0 1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_65
timestamp 0
transform 1 0 6532 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_77
timestamp 0
transform 1 0 7636 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_83
timestamp 0
transform 1 0 8188 0 1 12512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_85
timestamp 0
transform 1 0 8372 0 1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_97
timestamp 0
transform 1 0 9476 0 1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_109
timestamp 0
transform 1 0 10580 0 1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_121
timestamp 0
transform 1 0 11684 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_133
timestamp 0
transform 1 0 12788 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_139
timestamp 0
transform 1 0 13340 0 1 12512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_141
timestamp 0
transform 1 0 13524 0 1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_153
timestamp 0
transform 1 0 14628 0 1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_165
timestamp 0
transform 1 0 15732 0 1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_177
timestamp 0
transform 1 0 16836 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_189
timestamp 0
transform 1 0 17940 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_195
timestamp 0
transform 1 0 18492 0 1 12512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_197
timestamp 0
transform 1 0 18676 0 1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_209
timestamp 0
transform 1 0 19780 0 1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_221
timestamp 0
transform 1 0 20884 0 1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_233
timestamp 0
transform 1 0 21988 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_245
timestamp 0
transform 1 0 23092 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_251
timestamp 0
transform 1 0 23644 0 1 12512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_253
timestamp 0
transform 1 0 23828 0 1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_265
timestamp 0
transform 1 0 24932 0 1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_277
timestamp 0
transform 1 0 26036 0 1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_289
timestamp 0
transform 1 0 27140 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_301
timestamp 0
transform 1 0 28244 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_307
timestamp 0
transform 1 0 28796 0 1 12512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_309
timestamp 0
transform 1 0 28980 0 1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_321
timestamp 0
transform 1 0 30084 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_333
timestamp 0
transform 1 0 31188 0 1 12512
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_3
timestamp 0
transform 1 0 828 0 -1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_15
timestamp 0
transform 1 0 1932 0 -1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_27
timestamp 0
transform 1 0 3036 0 -1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_39
timestamp 0
transform 1 0 4140 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_51
timestamp 0
transform 1 0 5244 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_55
timestamp 0
transform 1 0 5612 0 -1 13600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_57
timestamp 0
transform 1 0 5796 0 -1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_69
timestamp 0
transform 1 0 6900 0 -1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_81
timestamp 0
transform 1 0 8004 0 -1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_93
timestamp 0
transform 1 0 9108 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_105
timestamp 0
transform 1 0 10212 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_111
timestamp 0
transform 1 0 10764 0 -1 13600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_113
timestamp 0
transform 1 0 10948 0 -1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_125
timestamp 0
transform 1 0 12052 0 -1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_137
timestamp 0
transform 1 0 13156 0 -1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_149
timestamp 0
transform 1 0 14260 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_161
timestamp 0
transform 1 0 15364 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_167
timestamp 0
transform 1 0 15916 0 -1 13600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_169
timestamp 0
transform 1 0 16100 0 -1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_181
timestamp 0
transform 1 0 17204 0 -1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_193
timestamp 0
transform 1 0 18308 0 -1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_205
timestamp 0
transform 1 0 19412 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_217
timestamp 0
transform 1 0 20516 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_223
timestamp 0
transform 1 0 21068 0 -1 13600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_225
timestamp 0
transform 1 0 21252 0 -1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_237
timestamp 0
transform 1 0 22356 0 -1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_249
timestamp 0
transform 1 0 23460 0 -1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_261
timestamp 0
transform 1 0 24564 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_273
timestamp 0
transform 1 0 25668 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_279
timestamp 0
transform 1 0 26220 0 -1 13600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_281
timestamp 0
transform 1 0 26404 0 -1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_293
timestamp 0
transform 1 0 27508 0 -1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_305
timestamp 0
transform 1 0 28612 0 -1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_317
timestamp 0
transform 1 0 29716 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_329
timestamp 0
transform 1 0 30820 0 -1 13600
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_3
timestamp 0
transform 1 0 828 0 1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_15
timestamp 0
transform 1 0 1932 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_27
timestamp 0
transform 1 0 3036 0 1 13600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_29
timestamp 0
transform 1 0 3220 0 1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_41
timestamp 0
transform 1 0 4324 0 1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_53
timestamp 0
transform 1 0 5428 0 1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_65
timestamp 0
transform 1 0 6532 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_77
timestamp 0
transform 1 0 7636 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_83
timestamp 0
transform 1 0 8188 0 1 13600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_85
timestamp 0
transform 1 0 8372 0 1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_97
timestamp 0
transform 1 0 9476 0 1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_109
timestamp 0
transform 1 0 10580 0 1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_121
timestamp 0
transform 1 0 11684 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_133
timestamp 0
transform 1 0 12788 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_139
timestamp 0
transform 1 0 13340 0 1 13600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_141
timestamp 0
transform 1 0 13524 0 1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_153
timestamp 0
transform 1 0 14628 0 1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_165
timestamp 0
transform 1 0 15732 0 1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_177
timestamp 0
transform 1 0 16836 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_189
timestamp 0
transform 1 0 17940 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_195
timestamp 0
transform 1 0 18492 0 1 13600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_197
timestamp 0
transform 1 0 18676 0 1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_209
timestamp 0
transform 1 0 19780 0 1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_221
timestamp 0
transform 1 0 20884 0 1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_233
timestamp 0
transform 1 0 21988 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_245
timestamp 0
transform 1 0 23092 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_251
timestamp 0
transform 1 0 23644 0 1 13600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_253
timestamp 0
transform 1 0 23828 0 1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_265
timestamp 0
transform 1 0 24932 0 1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_277
timestamp 0
transform 1 0 26036 0 1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_289
timestamp 0
transform 1 0 27140 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_301
timestamp 0
transform 1 0 28244 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_307
timestamp 0
transform 1 0 28796 0 1 13600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_309
timestamp 0
transform 1 0 28980 0 1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_321
timestamp 0
transform 1 0 30084 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_333
timestamp 0
transform 1 0 31188 0 1 13600
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_3
timestamp 0
transform 1 0 828 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_15
timestamp 0
transform 1 0 1932 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_27
timestamp 0
transform 1 0 3036 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_39
timestamp 0
transform 1 0 4140 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_51
timestamp 0
transform 1 0 5244 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_55
timestamp 0
transform 1 0 5612 0 -1 14688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_57
timestamp 0
transform 1 0 5796 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_69
timestamp 0
transform 1 0 6900 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_81
timestamp 0
transform 1 0 8004 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_93
timestamp 0
transform 1 0 9108 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_105
timestamp 0
transform 1 0 10212 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_111
timestamp 0
transform 1 0 10764 0 -1 14688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_113
timestamp 0
transform 1 0 10948 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_125
timestamp 0
transform 1 0 12052 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_137
timestamp 0
transform 1 0 13156 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_149
timestamp 0
transform 1 0 14260 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_161
timestamp 0
transform 1 0 15364 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_167
timestamp 0
transform 1 0 15916 0 -1 14688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_169
timestamp 0
transform 1 0 16100 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_181
timestamp 0
transform 1 0 17204 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_193
timestamp 0
transform 1 0 18308 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_205
timestamp 0
transform 1 0 19412 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_217
timestamp 0
transform 1 0 20516 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_223
timestamp 0
transform 1 0 21068 0 -1 14688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_225
timestamp 0
transform 1 0 21252 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_237
timestamp 0
transform 1 0 22356 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_249
timestamp 0
transform 1 0 23460 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_261
timestamp 0
transform 1 0 24564 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_273
timestamp 0
transform 1 0 25668 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_279
timestamp 0
transform 1 0 26220 0 -1 14688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_281
timestamp 0
transform 1 0 26404 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_293
timestamp 0
transform 1 0 27508 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_305
timestamp 0
transform 1 0 28612 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_317
timestamp 0
transform 1 0 29716 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_329
timestamp 0
transform 1 0 30820 0 -1 14688
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_3
timestamp 0
transform 1 0 828 0 1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_15
timestamp 0
transform 1 0 1932 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_27
timestamp 0
transform 1 0 3036 0 1 14688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_29
timestamp 0
transform 1 0 3220 0 1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_41
timestamp 0
transform 1 0 4324 0 1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_53
timestamp 0
transform 1 0 5428 0 1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_65
timestamp 0
transform 1 0 6532 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_77
timestamp 0
transform 1 0 7636 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_83
timestamp 0
transform 1 0 8188 0 1 14688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_85
timestamp 0
transform 1 0 8372 0 1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_97
timestamp 0
transform 1 0 9476 0 1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_109
timestamp 0
transform 1 0 10580 0 1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_121
timestamp 0
transform 1 0 11684 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_133
timestamp 0
transform 1 0 12788 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_139
timestamp 0
transform 1 0 13340 0 1 14688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_141
timestamp 0
transform 1 0 13524 0 1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_153
timestamp 0
transform 1 0 14628 0 1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_165
timestamp 0
transform 1 0 15732 0 1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_177
timestamp 0
transform 1 0 16836 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_189
timestamp 0
transform 1 0 17940 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_195
timestamp 0
transform 1 0 18492 0 1 14688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_197
timestamp 0
transform 1 0 18676 0 1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_209
timestamp 0
transform 1 0 19780 0 1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_221
timestamp 0
transform 1 0 20884 0 1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_233
timestamp 0
transform 1 0 21988 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_245
timestamp 0
transform 1 0 23092 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_251
timestamp 0
transform 1 0 23644 0 1 14688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_253
timestamp 0
transform 1 0 23828 0 1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_265
timestamp 0
transform 1 0 24932 0 1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_277
timestamp 0
transform 1 0 26036 0 1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_289
timestamp 0
transform 1 0 27140 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_301
timestamp 0
transform 1 0 28244 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_307
timestamp 0
transform 1 0 28796 0 1 14688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_309
timestamp 0
transform 1 0 28980 0 1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_321
timestamp 0
transform 1 0 30084 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_333
timestamp 0
transform 1 0 31188 0 1 14688
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_3
timestamp 0
transform 1 0 828 0 -1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_15
timestamp 0
transform 1 0 1932 0 -1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_27
timestamp 0
transform 1 0 3036 0 -1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_39
timestamp 0
transform 1 0 4140 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_51
timestamp 0
transform 1 0 5244 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_55
timestamp 0
transform 1 0 5612 0 -1 15776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_57
timestamp 0
transform 1 0 5796 0 -1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_69
timestamp 0
transform 1 0 6900 0 -1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_81
timestamp 0
transform 1 0 8004 0 -1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_93
timestamp 0
transform 1 0 9108 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_105
timestamp 0
transform 1 0 10212 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_111
timestamp 0
transform 1 0 10764 0 -1 15776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_113
timestamp 0
transform 1 0 10948 0 -1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_125
timestamp 0
transform 1 0 12052 0 -1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_137
timestamp 0
transform 1 0 13156 0 -1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_149
timestamp 0
transform 1 0 14260 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_161
timestamp 0
transform 1 0 15364 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_167
timestamp 0
transform 1 0 15916 0 -1 15776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_169
timestamp 0
transform 1 0 16100 0 -1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_181
timestamp 0
transform 1 0 17204 0 -1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_193
timestamp 0
transform 1 0 18308 0 -1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_205
timestamp 0
transform 1 0 19412 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_217
timestamp 0
transform 1 0 20516 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_223
timestamp 0
transform 1 0 21068 0 -1 15776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_225
timestamp 0
transform 1 0 21252 0 -1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_237
timestamp 0
transform 1 0 22356 0 -1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_249
timestamp 0
transform 1 0 23460 0 -1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_261
timestamp 0
transform 1 0 24564 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_273
timestamp 0
transform 1 0 25668 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_279
timestamp 0
transform 1 0 26220 0 -1 15776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_281
timestamp 0
transform 1 0 26404 0 -1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_293
timestamp 0
transform 1 0 27508 0 -1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_305
timestamp 0
transform 1 0 28612 0 -1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_317
timestamp 0
transform 1 0 29716 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_329
timestamp 0
transform 1 0 30820 0 -1 15776
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_3
timestamp 0
transform 1 0 828 0 1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_15
timestamp 0
transform 1 0 1932 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_27
timestamp 0
transform 1 0 3036 0 1 15776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_29
timestamp 0
transform 1 0 3220 0 1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_41
timestamp 0
transform 1 0 4324 0 1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_53
timestamp 0
transform 1 0 5428 0 1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_65
timestamp 0
transform 1 0 6532 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_77
timestamp 0
transform 1 0 7636 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_83
timestamp 0
transform 1 0 8188 0 1 15776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_85
timestamp 0
transform 1 0 8372 0 1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_97
timestamp 0
transform 1 0 9476 0 1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_109
timestamp 0
transform 1 0 10580 0 1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_121
timestamp 0
transform 1 0 11684 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_133
timestamp 0
transform 1 0 12788 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_139
timestamp 0
transform 1 0 13340 0 1 15776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_141
timestamp 0
transform 1 0 13524 0 1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_153
timestamp 0
transform 1 0 14628 0 1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_165
timestamp 0
transform 1 0 15732 0 1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_177
timestamp 0
transform 1 0 16836 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_189
timestamp 0
transform 1 0 17940 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_195
timestamp 0
transform 1 0 18492 0 1 15776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_197
timestamp 0
transform 1 0 18676 0 1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_209
timestamp 0
transform 1 0 19780 0 1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_221
timestamp 0
transform 1 0 20884 0 1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_233
timestamp 0
transform 1 0 21988 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_245
timestamp 0
transform 1 0 23092 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_251
timestamp 0
transform 1 0 23644 0 1 15776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_253
timestamp 0
transform 1 0 23828 0 1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_265
timestamp 0
transform 1 0 24932 0 1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_277
timestamp 0
transform 1 0 26036 0 1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_289
timestamp 0
transform 1 0 27140 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_301
timestamp 0
transform 1 0 28244 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_307
timestamp 0
transform 1 0 28796 0 1 15776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_309
timestamp 0
transform 1 0 28980 0 1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_321
timestamp 0
transform 1 0 30084 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_333
timestamp 0
transform 1 0 31188 0 1 15776
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_3
timestamp 0
transform 1 0 828 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_15
timestamp 0
transform 1 0 1932 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_27
timestamp 0
transform 1 0 3036 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_39
timestamp 0
transform 1 0 4140 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_51
timestamp 0
transform 1 0 5244 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_55
timestamp 0
transform 1 0 5612 0 -1 16864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_57
timestamp 0
transform 1 0 5796 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_69
timestamp 0
transform 1 0 6900 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_81
timestamp 0
transform 1 0 8004 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_93
timestamp 0
transform 1 0 9108 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_105
timestamp 0
transform 1 0 10212 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_111
timestamp 0
transform 1 0 10764 0 -1 16864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_113
timestamp 0
transform 1 0 10948 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_125
timestamp 0
transform 1 0 12052 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_137
timestamp 0
transform 1 0 13156 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_149
timestamp 0
transform 1 0 14260 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_161
timestamp 0
transform 1 0 15364 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_167
timestamp 0
transform 1 0 15916 0 -1 16864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_169
timestamp 0
transform 1 0 16100 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_181
timestamp 0
transform 1 0 17204 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_193
timestamp 0
transform 1 0 18308 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_205
timestamp 0
transform 1 0 19412 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_217
timestamp 0
transform 1 0 20516 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_223
timestamp 0
transform 1 0 21068 0 -1 16864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_225
timestamp 0
transform 1 0 21252 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_237
timestamp 0
transform 1 0 22356 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_249
timestamp 0
transform 1 0 23460 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_261
timestamp 0
transform 1 0 24564 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_273
timestamp 0
transform 1 0 25668 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_279
timestamp 0
transform 1 0 26220 0 -1 16864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_281
timestamp 0
transform 1 0 26404 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_293
timestamp 0
transform 1 0 27508 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_305
timestamp 0
transform 1 0 28612 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_317
timestamp 0
transform 1 0 29716 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_329
timestamp 0
transform 1 0 30820 0 -1 16864
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_3
timestamp 0
transform 1 0 828 0 1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_15
timestamp 0
transform 1 0 1932 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_27
timestamp 0
transform 1 0 3036 0 1 16864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_29
timestamp 0
transform 1 0 3220 0 1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_41
timestamp 0
transform 1 0 4324 0 1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_53
timestamp 0
transform 1 0 5428 0 1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_65
timestamp 0
transform 1 0 6532 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_77
timestamp 0
transform 1 0 7636 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_83
timestamp 0
transform 1 0 8188 0 1 16864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_85
timestamp 0
transform 1 0 8372 0 1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_97
timestamp 0
transform 1 0 9476 0 1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_109
timestamp 0
transform 1 0 10580 0 1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_121
timestamp 0
transform 1 0 11684 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_133
timestamp 0
transform 1 0 12788 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_139
timestamp 0
transform 1 0 13340 0 1 16864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_141
timestamp 0
transform 1 0 13524 0 1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_153
timestamp 0
transform 1 0 14628 0 1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_165
timestamp 0
transform 1 0 15732 0 1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_177
timestamp 0
transform 1 0 16836 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_189
timestamp 0
transform 1 0 17940 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_195
timestamp 0
transform 1 0 18492 0 1 16864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_197
timestamp 0
transform 1 0 18676 0 1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_209
timestamp 0
transform 1 0 19780 0 1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_221
timestamp 0
transform 1 0 20884 0 1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_233
timestamp 0
transform 1 0 21988 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_245
timestamp 0
transform 1 0 23092 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_251
timestamp 0
transform 1 0 23644 0 1 16864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_253
timestamp 0
transform 1 0 23828 0 1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_265
timestamp 0
transform 1 0 24932 0 1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_277
timestamp 0
transform 1 0 26036 0 1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_289
timestamp 0
transform 1 0 27140 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_301
timestamp 0
transform 1 0 28244 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_307
timestamp 0
transform 1 0 28796 0 1 16864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_309
timestamp 0
transform 1 0 28980 0 1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_321
timestamp 0
transform 1 0 30084 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_333
timestamp 0
transform 1 0 31188 0 1 16864
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_3
timestamp 0
transform 1 0 828 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_15
timestamp 0
transform 1 0 1932 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_27
timestamp 0
transform 1 0 3036 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_39
timestamp 0
transform 1 0 4140 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_51
timestamp 0
transform 1 0 5244 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_55
timestamp 0
transform 1 0 5612 0 -1 17952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_57
timestamp 0
transform 1 0 5796 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_69
timestamp 0
transform 1 0 6900 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_81
timestamp 0
transform 1 0 8004 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_93
timestamp 0
transform 1 0 9108 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_105
timestamp 0
transform 1 0 10212 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_111
timestamp 0
transform 1 0 10764 0 -1 17952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_113
timestamp 0
transform 1 0 10948 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_125
timestamp 0
transform 1 0 12052 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_137
timestamp 0
transform 1 0 13156 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_149
timestamp 0
transform 1 0 14260 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_161
timestamp 0
transform 1 0 15364 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_167
timestamp 0
transform 1 0 15916 0 -1 17952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_169
timestamp 0
transform 1 0 16100 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_181
timestamp 0
transform 1 0 17204 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_193
timestamp 0
transform 1 0 18308 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_205
timestamp 0
transform 1 0 19412 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_217
timestamp 0
transform 1 0 20516 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_223
timestamp 0
transform 1 0 21068 0 -1 17952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_225
timestamp 0
transform 1 0 21252 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_237
timestamp 0
transform 1 0 22356 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_249
timestamp 0
transform 1 0 23460 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_261
timestamp 0
transform 1 0 24564 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_273
timestamp 0
transform 1 0 25668 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_279
timestamp 0
transform 1 0 26220 0 -1 17952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_281
timestamp 0
transform 1 0 26404 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_293
timestamp 0
transform 1 0 27508 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_305
timestamp 0
transform 1 0 28612 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_317
timestamp 0
transform 1 0 29716 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_329
timestamp 0
transform 1 0 30820 0 -1 17952
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_3
timestamp 0
transform 1 0 828 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_15
timestamp 0
transform 1 0 1932 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_27
timestamp 0
transform 1 0 3036 0 1 17952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_29
timestamp 0
transform 1 0 3220 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_41
timestamp 0
transform 1 0 4324 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_53
timestamp 0
transform 1 0 5428 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_65
timestamp 0
transform 1 0 6532 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_77
timestamp 0
transform 1 0 7636 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_83
timestamp 0
transform 1 0 8188 0 1 17952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_85
timestamp 0
transform 1 0 8372 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_97
timestamp 0
transform 1 0 9476 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_109
timestamp 0
transform 1 0 10580 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_121
timestamp 0
transform 1 0 11684 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_133
timestamp 0
transform 1 0 12788 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_139
timestamp 0
transform 1 0 13340 0 1 17952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_141
timestamp 0
transform 1 0 13524 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_153
timestamp 0
transform 1 0 14628 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_165
timestamp 0
transform 1 0 15732 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_177
timestamp 0
transform 1 0 16836 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_189
timestamp 0
transform 1 0 17940 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_195
timestamp 0
transform 1 0 18492 0 1 17952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_197
timestamp 0
transform 1 0 18676 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_209
timestamp 0
transform 1 0 19780 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_221
timestamp 0
transform 1 0 20884 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_233
timestamp 0
transform 1 0 21988 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_245
timestamp 0
transform 1 0 23092 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_251
timestamp 0
transform 1 0 23644 0 1 17952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_253
timestamp 0
transform 1 0 23828 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_265
timestamp 0
transform 1 0 24932 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_277
timestamp 0
transform 1 0 26036 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_289
timestamp 0
transform 1 0 27140 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_301
timestamp 0
transform 1 0 28244 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_307
timestamp 0
transform 1 0 28796 0 1 17952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_309
timestamp 0
transform 1 0 28980 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_321
timestamp 0
transform 1 0 30084 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_333
timestamp 0
transform 1 0 31188 0 1 17952
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_3
timestamp 0
transform 1 0 828 0 -1 19040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_15
timestamp 0
transform 1 0 1932 0 -1 19040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_27
timestamp 0
transform 1 0 3036 0 -1 19040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_39
timestamp 0
transform 1 0 4140 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_51
timestamp 0
transform 1 0 5244 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_55
timestamp 0
transform 1 0 5612 0 -1 19040
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_57
timestamp 0
transform 1 0 5796 0 -1 19040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_69
timestamp 0
transform 1 0 6900 0 -1 19040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_81
timestamp 0
transform 1 0 8004 0 -1 19040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_93
timestamp 0
transform 1 0 9108 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_105
timestamp 0
transform 1 0 10212 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_111
timestamp 0
transform 1 0 10764 0 -1 19040
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_113
timestamp 0
transform 1 0 10948 0 -1 19040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_125
timestamp 0
transform 1 0 12052 0 -1 19040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_137
timestamp 0
transform 1 0 13156 0 -1 19040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_149
timestamp 0
transform 1 0 14260 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_161
timestamp 0
transform 1 0 15364 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_167
timestamp 0
transform 1 0 15916 0 -1 19040
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_169
timestamp 0
transform 1 0 16100 0 -1 19040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_181
timestamp 0
transform 1 0 17204 0 -1 19040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_193
timestamp 0
transform 1 0 18308 0 -1 19040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_205
timestamp 0
transform 1 0 19412 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_217
timestamp 0
transform 1 0 20516 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_223
timestamp 0
transform 1 0 21068 0 -1 19040
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_225
timestamp 0
transform 1 0 21252 0 -1 19040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_237
timestamp 0
transform 1 0 22356 0 -1 19040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_249
timestamp 0
transform 1 0 23460 0 -1 19040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_261
timestamp 0
transform 1 0 24564 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_273
timestamp 0
transform 1 0 25668 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_279
timestamp 0
transform 1 0 26220 0 -1 19040
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_281
timestamp 0
transform 1 0 26404 0 -1 19040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_293
timestamp 0
transform 1 0 27508 0 -1 19040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_305
timestamp 0
transform 1 0 28612 0 -1 19040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_317
timestamp 0
transform 1 0 29716 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_329
timestamp 0
transform 1 0 30820 0 -1 19040
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_3
timestamp 0
transform 1 0 828 0 1 19040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_15
timestamp 0
transform 1 0 1932 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_27
timestamp 0
transform 1 0 3036 0 1 19040
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_29
timestamp 0
transform 1 0 3220 0 1 19040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_41
timestamp 0
transform 1 0 4324 0 1 19040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_53
timestamp 0
transform 1 0 5428 0 1 19040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_65
timestamp 0
transform 1 0 6532 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_77
timestamp 0
transform 1 0 7636 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_83
timestamp 0
transform 1 0 8188 0 1 19040
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_85
timestamp 0
transform 1 0 8372 0 1 19040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_97
timestamp 0
transform 1 0 9476 0 1 19040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_109
timestamp 0
transform 1 0 10580 0 1 19040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_121
timestamp 0
transform 1 0 11684 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_133
timestamp 0
transform 1 0 12788 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_139
timestamp 0
transform 1 0 13340 0 1 19040
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_141
timestamp 0
transform 1 0 13524 0 1 19040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_153
timestamp 0
transform 1 0 14628 0 1 19040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_165
timestamp 0
transform 1 0 15732 0 1 19040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_177
timestamp 0
transform 1 0 16836 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_189
timestamp 0
transform 1 0 17940 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_195
timestamp 0
transform 1 0 18492 0 1 19040
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_197
timestamp 0
transform 1 0 18676 0 1 19040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_209
timestamp 0
transform 1 0 19780 0 1 19040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_221
timestamp 0
transform 1 0 20884 0 1 19040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_233
timestamp 0
transform 1 0 21988 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_245
timestamp 0
transform 1 0 23092 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_251
timestamp 0
transform 1 0 23644 0 1 19040
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_253
timestamp 0
transform 1 0 23828 0 1 19040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_265
timestamp 0
transform 1 0 24932 0 1 19040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_277
timestamp 0
transform 1 0 26036 0 1 19040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_289
timestamp 0
transform 1 0 27140 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_301
timestamp 0
transform 1 0 28244 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_307
timestamp 0
transform 1 0 28796 0 1 19040
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_309
timestamp 0
transform 1 0 28980 0 1 19040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_321
timestamp 0
transform 1 0 30084 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_333
timestamp 0
transform 1 0 31188 0 1 19040
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_3
timestamp 0
transform 1 0 828 0 -1 20128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_15
timestamp 0
transform 1 0 1932 0 -1 20128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_27
timestamp 0
transform 1 0 3036 0 -1 20128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_39
timestamp 0
transform 1 0 4140 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_51
timestamp 0
transform 1 0 5244 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_55
timestamp 0
transform 1 0 5612 0 -1 20128
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_57
timestamp 0
transform 1 0 5796 0 -1 20128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_69
timestamp 0
transform 1 0 6900 0 -1 20128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_81
timestamp 0
transform 1 0 8004 0 -1 20128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_93
timestamp 0
transform 1 0 9108 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_105
timestamp 0
transform 1 0 10212 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_111
timestamp 0
transform 1 0 10764 0 -1 20128
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_113
timestamp 0
transform 1 0 10948 0 -1 20128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_125
timestamp 0
transform 1 0 12052 0 -1 20128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_137
timestamp 0
transform 1 0 13156 0 -1 20128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_149
timestamp 0
transform 1 0 14260 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_161
timestamp 0
transform 1 0 15364 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_167
timestamp 0
transform 1 0 15916 0 -1 20128
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_169
timestamp 0
transform 1 0 16100 0 -1 20128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_181
timestamp 0
transform 1 0 17204 0 -1 20128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_193
timestamp 0
transform 1 0 18308 0 -1 20128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_205
timestamp 0
transform 1 0 19412 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_217
timestamp 0
transform 1 0 20516 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_223
timestamp 0
transform 1 0 21068 0 -1 20128
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_225
timestamp 0
transform 1 0 21252 0 -1 20128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_237
timestamp 0
transform 1 0 22356 0 -1 20128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_249
timestamp 0
transform 1 0 23460 0 -1 20128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_261
timestamp 0
transform 1 0 24564 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_273
timestamp 0
transform 1 0 25668 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_279
timestamp 0
transform 1 0 26220 0 -1 20128
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_281
timestamp 0
transform 1 0 26404 0 -1 20128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_293
timestamp 0
transform 1 0 27508 0 -1 20128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_305
timestamp 0
transform 1 0 28612 0 -1 20128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_317
timestamp 0
transform 1 0 29716 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_329
timestamp 0
transform 1 0 30820 0 -1 20128
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_3
timestamp 0
transform 1 0 828 0 1 20128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_15
timestamp 0
transform 1 0 1932 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_27
timestamp 0
transform 1 0 3036 0 1 20128
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_29
timestamp 0
transform 1 0 3220 0 1 20128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_41
timestamp 0
transform 1 0 4324 0 1 20128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_53
timestamp 0
transform 1 0 5428 0 1 20128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_65
timestamp 0
transform 1 0 6532 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_77
timestamp 0
transform 1 0 7636 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_83
timestamp 0
transform 1 0 8188 0 1 20128
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_85
timestamp 0
transform 1 0 8372 0 1 20128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_97
timestamp 0
transform 1 0 9476 0 1 20128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_109
timestamp 0
transform 1 0 10580 0 1 20128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_121
timestamp 0
transform 1 0 11684 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_133
timestamp 0
transform 1 0 12788 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_139
timestamp 0
transform 1 0 13340 0 1 20128
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_141
timestamp 0
transform 1 0 13524 0 1 20128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_153
timestamp 0
transform 1 0 14628 0 1 20128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_165
timestamp 0
transform 1 0 15732 0 1 20128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_177
timestamp 0
transform 1 0 16836 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_189
timestamp 0
transform 1 0 17940 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_195
timestamp 0
transform 1 0 18492 0 1 20128
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_197
timestamp 0
transform 1 0 18676 0 1 20128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_209
timestamp 0
transform 1 0 19780 0 1 20128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_221
timestamp 0
transform 1 0 20884 0 1 20128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_233
timestamp 0
transform 1 0 21988 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_245
timestamp 0
transform 1 0 23092 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_251
timestamp 0
transform 1 0 23644 0 1 20128
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_253
timestamp 0
transform 1 0 23828 0 1 20128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_265
timestamp 0
transform 1 0 24932 0 1 20128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_277
timestamp 0
transform 1 0 26036 0 1 20128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_289
timestamp 0
transform 1 0 27140 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_301
timestamp 0
transform 1 0 28244 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_307
timestamp 0
transform 1 0 28796 0 1 20128
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_309
timestamp 0
transform 1 0 28980 0 1 20128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_321
timestamp 0
transform 1 0 30084 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_333
timestamp 0
transform 1 0 31188 0 1 20128
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_3
timestamp 0
transform 1 0 828 0 -1 21216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_15
timestamp 0
transform 1 0 1932 0 -1 21216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_27
timestamp 0
transform 1 0 3036 0 -1 21216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_39
timestamp 0
transform 1 0 4140 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_51
timestamp 0
transform 1 0 5244 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_55
timestamp 0
transform 1 0 5612 0 -1 21216
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_57
timestamp 0
transform 1 0 5796 0 -1 21216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_69
timestamp 0
transform 1 0 6900 0 -1 21216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_81
timestamp 0
transform 1 0 8004 0 -1 21216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_93
timestamp 0
transform 1 0 9108 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_105
timestamp 0
transform 1 0 10212 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_111
timestamp 0
transform 1 0 10764 0 -1 21216
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_113
timestamp 0
transform 1 0 10948 0 -1 21216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_125
timestamp 0
transform 1 0 12052 0 -1 21216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_137
timestamp 0
transform 1 0 13156 0 -1 21216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_149
timestamp 0
transform 1 0 14260 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_161
timestamp 0
transform 1 0 15364 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_167
timestamp 0
transform 1 0 15916 0 -1 21216
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_169
timestamp 0
transform 1 0 16100 0 -1 21216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_181
timestamp 0
transform 1 0 17204 0 -1 21216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_193
timestamp 0
transform 1 0 18308 0 -1 21216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_205
timestamp 0
transform 1 0 19412 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_217
timestamp 0
transform 1 0 20516 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_223
timestamp 0
transform 1 0 21068 0 -1 21216
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_225
timestamp 0
transform 1 0 21252 0 -1 21216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_237
timestamp 0
transform 1 0 22356 0 -1 21216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_249
timestamp 0
transform 1 0 23460 0 -1 21216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_261
timestamp 0
transform 1 0 24564 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_273
timestamp 0
transform 1 0 25668 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_279
timestamp 0
transform 1 0 26220 0 -1 21216
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_281
timestamp 0
transform 1 0 26404 0 -1 21216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_293
timestamp 0
transform 1 0 27508 0 -1 21216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_305
timestamp 0
transform 1 0 28612 0 -1 21216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_317
timestamp 0
transform 1 0 29716 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_329
timestamp 0
transform 1 0 30820 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_6
timestamp 0
transform 1 0 1104 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_10
timestamp 0
transform 1 0 1472 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_14
timestamp 0
transform 1 0 1840 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_18
timestamp 0
transform 1 0 2208 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_22
timestamp 0
transform 1 0 2576 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_32
timestamp 0
transform 1 0 3496 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_38
timestamp 0
transform 1 0 4048 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_42
timestamp 0
transform 1 0 4416 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_46
timestamp 0
transform 1 0 4784 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_50
timestamp 0
transform 1 0 5152 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_54
timestamp 0
transform 1 0 5520 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_57
timestamp 0
transform 1 0 5796 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_62
timestamp 0
transform 1 0 6256 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_66
timestamp 0
transform 1 0 6624 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_70
timestamp 0
transform 1 0 6992 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_74
timestamp 0
transform 1 0 7360 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_78
timestamp 0
transform 1 0 7728 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_88
timestamp 0
transform 1 0 8648 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_94
timestamp 0
transform 1 0 9200 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_98
timestamp 0
transform 1 0 9568 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_102
timestamp 0
transform 1 0 9936 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_106
timestamp 0
transform 1 0 10304 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_110
timestamp 0
transform 1 0 10672 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_113
timestamp 0
transform 1 0 10948 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_118
timestamp 0
transform 1 0 11408 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_122
timestamp 0
transform 1 0 11776 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_126
timestamp 0
transform 1 0 12144 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_130
timestamp 0
transform 1 0 12512 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_134
timestamp 0
transform 1 0 12880 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_144
timestamp 0
transform 1 0 13800 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_150
timestamp 0
transform 1 0 14352 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_154
timestamp 0
transform 1 0 14720 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_158
timestamp 0
transform 1 0 15088 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_162
timestamp 0
transform 1 0 15456 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_166
timestamp 0
transform 1 0 15824 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_169
timestamp 0
transform 1 0 16100 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_174
timestamp 0
transform 1 0 16560 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_178
timestamp 0
transform 1 0 16928 0 1 21216
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_182
timestamp 0
transform 1 0 17296 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_194
timestamp 0
transform 1 0 18400 0 1 21216
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_197
timestamp 0
transform 1 0 18676 0 1 21216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_209
timestamp 0
transform 1 0 19780 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_221
timestamp 0
transform 1 0 20884 0 1 21216
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_225
timestamp 0
transform 1 0 21252 0 1 21216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_237
timestamp 0
transform 1 0 22356 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_249
timestamp 0
transform 1 0 23460 0 1 21216
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_253
timestamp 0
transform 1 0 23828 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_265
timestamp 0
transform 1 0 24932 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_271
timestamp 0
transform 1 0 25484 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_278
timestamp 0
transform 1 0 26128 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_281
timestamp 0
transform 1 0 26404 0 1 21216
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_290
timestamp 0
transform 1 0 27232 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_302
timestamp 0
transform 1 0 28336 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_312
timestamp 0
transform 1 0 29256 0 1 21216
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_318
timestamp 0
transform 1 0 29808 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_330
timestamp 0
transform 1 0 30912 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_334
timestamp 0
transform 1 0 31280 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 0
transform 1 0 29532 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 0
transform 1 0 28980 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_39
timestamp 0
transform 1 0 552 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 0
transform -1 0 31648 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_40
timestamp 0
transform 1 0 552 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 0
transform -1 0 31648 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_41
timestamp 0
transform 1 0 552 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 0
transform -1 0 31648 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_42
timestamp 0
transform 1 0 552 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp 0
transform -1 0 31648 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_43
timestamp 0
transform 1 0 552 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp 0
transform -1 0 31648 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_44
timestamp 0
transform 1 0 552 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp 0
transform -1 0 31648 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_45
timestamp 0
transform 1 0 552 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp 0
transform -1 0 31648 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_46
timestamp 0
transform 1 0 552 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp 0
transform -1 0 31648 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_47
timestamp 0
transform 1 0 552 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp 0
transform -1 0 31648 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_48
timestamp 0
transform 1 0 552 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp 0
transform -1 0 31648 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_49
timestamp 0
transform 1 0 552 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp 0
transform -1 0 31648 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_50
timestamp 0
transform 1 0 552 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp 0
transform -1 0 31648 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Left_51
timestamp 0
transform 1 0 552 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Right_12
timestamp 0
transform -1 0 31648 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Left_52
timestamp 0
transform 1 0 552 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Right_13
timestamp 0
transform -1 0 31648 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Left_53
timestamp 0
transform 1 0 552 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Right_14
timestamp 0
transform -1 0 31648 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Left_54
timestamp 0
transform 1 0 552 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Right_15
timestamp 0
transform -1 0 31648 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Left_55
timestamp 0
transform 1 0 552 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Right_16
timestamp 0
transform -1 0 31648 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Left_56
timestamp 0
transform 1 0 552 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Right_17
timestamp 0
transform -1 0 31648 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Left_57
timestamp 0
transform 1 0 552 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Right_18
timestamp 0
transform -1 0 31648 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Left_58
timestamp 0
transform 1 0 552 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Right_19
timestamp 0
transform -1 0 31648 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Left_59
timestamp 0
transform 1 0 552 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Right_20
timestamp 0
transform -1 0 31648 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Left_60
timestamp 0
transform 1 0 552 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Right_21
timestamp 0
transform -1 0 31648 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Left_61
timestamp 0
transform 1 0 552 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Right_22
timestamp 0
transform -1 0 31648 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Left_62
timestamp 0
transform 1 0 552 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Right_23
timestamp 0
transform -1 0 31648 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Left_63
timestamp 0
transform 1 0 552 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Right_24
timestamp 0
transform -1 0 31648 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Left_64
timestamp 0
transform 1 0 552 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Right_25
timestamp 0
transform -1 0 31648 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Left_65
timestamp 0
transform 1 0 552 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Right_26
timestamp 0
transform -1 0 31648 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Left_66
timestamp 0
transform 1 0 552 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Right_27
timestamp 0
transform -1 0 31648 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Left_67
timestamp 0
transform 1 0 552 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Right_28
timestamp 0
transform -1 0 31648 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Left_68
timestamp 0
transform 1 0 552 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Right_29
timestamp 0
transform -1 0 31648 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Left_69
timestamp 0
transform 1 0 552 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Right_30
timestamp 0
transform -1 0 31648 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_Left_70
timestamp 0
transform 1 0 552 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_Right_31
timestamp 0
transform -1 0 31648 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_Left_71
timestamp 0
transform 1 0 552 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_Right_32
timestamp 0
transform -1 0 31648 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_Left_72
timestamp 0
transform 1 0 552 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_Right_33
timestamp 0
transform -1 0 31648 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_Left_73
timestamp 0
transform 1 0 552 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_Right_34
timestamp 0
transform -1 0 31648 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_Left_74
timestamp 0
transform 1 0 552 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_Right_35
timestamp 0
transform -1 0 31648 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_Left_75
timestamp 0
transform 1 0 552 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_Right_36
timestamp 0
transform -1 0 31648 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_Left_76
timestamp 0
transform 1 0 552 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_Right_37
timestamp 0
transform -1 0 31648 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_Left_77
timestamp 0
transform 1 0 552 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_Right_38
timestamp 0
transform -1 0 31648 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_78
timestamp 0
transform 1 0 3128 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_79
timestamp 0
transform 1 0 5704 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_80
timestamp 0
transform 1 0 8280 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_81
timestamp 0
transform 1 0 10856 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_82
timestamp 0
transform 1 0 13432 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_83
timestamp 0
transform 1 0 16008 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_84
timestamp 0
transform 1 0 18584 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_85
timestamp 0
transform 1 0 21160 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_86
timestamp 0
transform 1 0 23736 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_87
timestamp 0
transform 1 0 26312 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_88
timestamp 0
transform 1 0 28888 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_89
timestamp 0
transform 1 0 5704 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_90
timestamp 0
transform 1 0 10856 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_91
timestamp 0
transform 1 0 16008 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_92
timestamp 0
transform 1 0 21160 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_93
timestamp 0
transform 1 0 26312 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_94
timestamp 0
transform 1 0 3128 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_95
timestamp 0
transform 1 0 8280 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_96
timestamp 0
transform 1 0 13432 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_97
timestamp 0
transform 1 0 18584 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_98
timestamp 0
transform 1 0 23736 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_99
timestamp 0
transform 1 0 28888 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_100
timestamp 0
transform 1 0 5704 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_101
timestamp 0
transform 1 0 10856 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_102
timestamp 0
transform 1 0 16008 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_103
timestamp 0
transform 1 0 21160 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_104
timestamp 0
transform 1 0 26312 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_105
timestamp 0
transform 1 0 3128 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_106
timestamp 0
transform 1 0 8280 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_107
timestamp 0
transform 1 0 13432 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_108
timestamp 0
transform 1 0 18584 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_109
timestamp 0
transform 1 0 23736 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_110
timestamp 0
transform 1 0 28888 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_111
timestamp 0
transform 1 0 5704 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_112
timestamp 0
transform 1 0 10856 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_113
timestamp 0
transform 1 0 16008 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_114
timestamp 0
transform 1 0 21160 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_115
timestamp 0
transform 1 0 26312 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_116
timestamp 0
transform 1 0 3128 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_117
timestamp 0
transform 1 0 8280 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_118
timestamp 0
transform 1 0 13432 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_119
timestamp 0
transform 1 0 18584 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_120
timestamp 0
transform 1 0 23736 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_121
timestamp 0
transform 1 0 28888 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_122
timestamp 0
transform 1 0 5704 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_123
timestamp 0
transform 1 0 10856 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_124
timestamp 0
transform 1 0 16008 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_125
timestamp 0
transform 1 0 21160 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_126
timestamp 0
transform 1 0 26312 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_127
timestamp 0
transform 1 0 3128 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_128
timestamp 0
transform 1 0 8280 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_129
timestamp 0
transform 1 0 13432 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_130
timestamp 0
transform 1 0 18584 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_131
timestamp 0
transform 1 0 23736 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_132
timestamp 0
transform 1 0 28888 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_133
timestamp 0
transform 1 0 5704 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_134
timestamp 0
transform 1 0 10856 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_135
timestamp 0
transform 1 0 16008 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_136
timestamp 0
transform 1 0 21160 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_137
timestamp 0
transform 1 0 26312 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_138
timestamp 0
transform 1 0 3128 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_139
timestamp 0
transform 1 0 8280 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_140
timestamp 0
transform 1 0 13432 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_141
timestamp 0
transform 1 0 18584 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_142
timestamp 0
transform 1 0 23736 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_143
timestamp 0
transform 1 0 28888 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_144
timestamp 0
transform 1 0 5704 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_145
timestamp 0
transform 1 0 10856 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_146
timestamp 0
transform 1 0 16008 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_147
timestamp 0
transform 1 0 21160 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_148
timestamp 0
transform 1 0 26312 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_149
timestamp 0
transform 1 0 3128 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_150
timestamp 0
transform 1 0 8280 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_151
timestamp 0
transform 1 0 13432 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_152
timestamp 0
transform 1 0 18584 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_153
timestamp 0
transform 1 0 23736 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_154
timestamp 0
transform 1 0 28888 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_155
timestamp 0
transform 1 0 5704 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_156
timestamp 0
transform 1 0 10856 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_157
timestamp 0
transform 1 0 16008 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_158
timestamp 0
transform 1 0 21160 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_159
timestamp 0
transform 1 0 26312 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_160
timestamp 0
transform 1 0 3128 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_161
timestamp 0
transform 1 0 8280 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_162
timestamp 0
transform 1 0 13432 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_163
timestamp 0
transform 1 0 18584 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_164
timestamp 0
transform 1 0 23736 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_165
timestamp 0
transform 1 0 28888 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_166
timestamp 0
transform 1 0 5704 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_167
timestamp 0
transform 1 0 10856 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_168
timestamp 0
transform 1 0 16008 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_169
timestamp 0
transform 1 0 21160 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_170
timestamp 0
transform 1 0 26312 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_171
timestamp 0
transform 1 0 3128 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_172
timestamp 0
transform 1 0 8280 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_173
timestamp 0
transform 1 0 13432 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_174
timestamp 0
transform 1 0 18584 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_175
timestamp 0
transform 1 0 23736 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_176
timestamp 0
transform 1 0 28888 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_177
timestamp 0
transform 1 0 5704 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_178
timestamp 0
transform 1 0 10856 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_179
timestamp 0
transform 1 0 16008 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_180
timestamp 0
transform 1 0 21160 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_181
timestamp 0
transform 1 0 26312 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_182
timestamp 0
transform 1 0 3128 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_183
timestamp 0
transform 1 0 8280 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_184
timestamp 0
transform 1 0 13432 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_185
timestamp 0
transform 1 0 18584 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_186
timestamp 0
transform 1 0 23736 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_187
timestamp 0
transform 1 0 28888 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_188
timestamp 0
transform 1 0 5704 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_189
timestamp 0
transform 1 0 10856 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_190
timestamp 0
transform 1 0 16008 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_191
timestamp 0
transform 1 0 21160 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_192
timestamp 0
transform 1 0 26312 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_193
timestamp 0
transform 1 0 3128 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_194
timestamp 0
transform 1 0 8280 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_195
timestamp 0
transform 1 0 13432 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_196
timestamp 0
transform 1 0 18584 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_197
timestamp 0
transform 1 0 23736 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_198
timestamp 0
transform 1 0 28888 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_199
timestamp 0
transform 1 0 5704 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_200
timestamp 0
transform 1 0 10856 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_201
timestamp 0
transform 1 0 16008 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_202
timestamp 0
transform 1 0 21160 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_203
timestamp 0
transform 1 0 26312 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_204
timestamp 0
transform 1 0 3128 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_205
timestamp 0
transform 1 0 8280 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_206
timestamp 0
transform 1 0 13432 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_207
timestamp 0
transform 1 0 18584 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_208
timestamp 0
transform 1 0 23736 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_209
timestamp 0
transform 1 0 28888 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_210
timestamp 0
transform 1 0 5704 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_211
timestamp 0
transform 1 0 10856 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_212
timestamp 0
transform 1 0 16008 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_213
timestamp 0
transform 1 0 21160 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_214
timestamp 0
transform 1 0 26312 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_215
timestamp 0
transform 1 0 3128 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_216
timestamp 0
transform 1 0 8280 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_217
timestamp 0
transform 1 0 13432 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_218
timestamp 0
transform 1 0 18584 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_219
timestamp 0
transform 1 0 23736 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_220
timestamp 0
transform 1 0 28888 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_221
timestamp 0
transform 1 0 5704 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_222
timestamp 0
transform 1 0 10856 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_223
timestamp 0
transform 1 0 16008 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_224
timestamp 0
transform 1 0 21160 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_225
timestamp 0
transform 1 0 26312 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_226
timestamp 0
transform 1 0 3128 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_227
timestamp 0
transform 1 0 8280 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_228
timestamp 0
transform 1 0 13432 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_229
timestamp 0
transform 1 0 18584 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_230
timestamp 0
transform 1 0 23736 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_231
timestamp 0
transform 1 0 28888 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_232
timestamp 0
transform 1 0 5704 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_233
timestamp 0
transform 1 0 10856 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_234
timestamp 0
transform 1 0 16008 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_235
timestamp 0
transform 1 0 21160 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_236
timestamp 0
transform 1 0 26312 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_237
timestamp 0
transform 1 0 3128 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_238
timestamp 0
transform 1 0 8280 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_239
timestamp 0
transform 1 0 13432 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_240
timestamp 0
transform 1 0 18584 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_241
timestamp 0
transform 1 0 23736 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_242
timestamp 0
transform 1 0 28888 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_243
timestamp 0
transform 1 0 5704 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_244
timestamp 0
transform 1 0 10856 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_245
timestamp 0
transform 1 0 16008 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_246
timestamp 0
transform 1 0 21160 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_247
timestamp 0
transform 1 0 26312 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_248
timestamp 0
transform 1 0 3128 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_249
timestamp 0
transform 1 0 8280 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_250
timestamp 0
transform 1 0 13432 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_251
timestamp 0
transform 1 0 18584 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_252
timestamp 0
transform 1 0 23736 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_253
timestamp 0
transform 1 0 28888 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_254
timestamp 0
transform 1 0 5704 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_255
timestamp 0
transform 1 0 10856 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_256
timestamp 0
transform 1 0 16008 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_257
timestamp 0
transform 1 0 21160 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_258
timestamp 0
transform 1 0 26312 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_259
timestamp 0
transform 1 0 3128 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_260
timestamp 0
transform 1 0 8280 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_261
timestamp 0
transform 1 0 13432 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_262
timestamp 0
transform 1 0 18584 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_263
timestamp 0
transform 1 0 23736 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_264
timestamp 0
transform 1 0 28888 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_265
timestamp 0
transform 1 0 5704 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_266
timestamp 0
transform 1 0 10856 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_267
timestamp 0
transform 1 0 16008 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_268
timestamp 0
transform 1 0 21160 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_269
timestamp 0
transform 1 0 26312 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_270
timestamp 0
transform 1 0 3128 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_271
timestamp 0
transform 1 0 8280 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_272
timestamp 0
transform 1 0 13432 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_273
timestamp 0
transform 1 0 18584 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_274
timestamp 0
transform 1 0 23736 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_275
timestamp 0
transform 1 0 28888 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_276
timestamp 0
transform 1 0 5704 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_277
timestamp 0
transform 1 0 10856 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_278
timestamp 0
transform 1 0 16008 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_279
timestamp 0
transform 1 0 21160 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_280
timestamp 0
transform 1 0 26312 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_281
timestamp 0
transform 1 0 3128 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_282
timestamp 0
transform 1 0 8280 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_283
timestamp 0
transform 1 0 13432 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_284
timestamp 0
transform 1 0 18584 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_285
timestamp 0
transform 1 0 23736 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_286
timestamp 0
transform 1 0 28888 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_287
timestamp 0
transform 1 0 5704 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_288
timestamp 0
transform 1 0 10856 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_289
timestamp 0
transform 1 0 16008 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_290
timestamp 0
transform 1 0 21160 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_291
timestamp 0
transform 1 0 26312 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_292
timestamp 0
transform 1 0 3128 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_293
timestamp 0
transform 1 0 5704 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_294
timestamp 0
transform 1 0 8280 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_295
timestamp 0
transform 1 0 10856 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_296
timestamp 0
transform 1 0 13432 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_297
timestamp 0
transform 1 0 16008 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_298
timestamp 0
transform 1 0 18584 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_299
timestamp 0
transform 1 0 21160 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_300
timestamp 0
transform 1 0 23736 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_301
timestamp 0
transform 1 0 26312 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_302
timestamp 0
transform 1 0 28888 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  tt_um_example_3
timestamp 0
transform -1 0 1104 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_example_4
timestamp 0
transform -1 0 12144 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_example_5
timestamp 0
transform -1 0 11408 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_example_6
timestamp 0
transform -1 0 10672 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_example_7
timestamp 0
transform -1 0 9936 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_example_8
timestamp 0
transform -1 0 9200 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_example_9
timestamp 0
transform -1 0 8648 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_example_10
timestamp 0
transform -1 0 7728 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_example_11
timestamp 0
transform -1 0 6992 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_example_12
timestamp 0
transform -1 0 17296 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_example_13
timestamp 0
transform -1 0 16560 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_example_14
timestamp 0
transform -1 0 15824 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_example_15
timestamp 0
transform -1 0 15088 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_example_16
timestamp 0
transform -1 0 14352 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_example_17
timestamp 0
transform -1 0 13800 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_example_18
timestamp 0
transform -1 0 12880 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_example_19
timestamp 0
transform -1 0 6256 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_example_20
timestamp 0
transform -1 0 5520 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_example_21
timestamp 0
transform -1 0 4784 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_example_22
timestamp 0
transform -1 0 4048 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_example_23
timestamp 0
transform -1 0 3496 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_example_24
timestamp 0
transform -1 0 2576 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_example_25
timestamp 0
transform -1 0 1840 0 1 21216
box -38 -48 314 592
<< labels >>
rlabel metal2 s 16180 21216 16180 21216 4 VGND
rlabel metal1 s 16100 21760 16100 21760 4 VPWR
rlabel metal1 s 26404 21386 26404 21386 4 _00_
rlabel metal2 s 27002 21658 27002 21658 4 net1
rlabel metal2 s 7498 21743 7498 21743 4 net10
rlabel metal2 s 6762 21743 6762 21743 4 net11
rlabel metal2 s 17066 21743 17066 21743 4 net12
rlabel metal2 s 16330 21811 16330 21811 4 net13
rlabel metal2 s 15594 21743 15594 21743 4 net14
rlabel metal2 s 14858 21743 14858 21743 4 net15
rlabel metal2 s 14122 21743 14122 21743 4 net16
rlabel metal2 s 13570 21743 13570 21743 4 net17
rlabel metal2 s 12650 21743 12650 21743 4 net18
rlabel metal2 s 6026 21743 6026 21743 4 net19
rlabel metal2 s 27186 21726 27186 21726 4 net2
rlabel metal2 s 5290 21743 5290 21743 4 net20
rlabel metal1 s 4600 21658 4600 21658 4 net21
rlabel metal2 s 3818 21743 3818 21743 4 net22
rlabel metal2 s 3266 21743 3266 21743 4 net23
rlabel metal2 s 2346 21743 2346 21743 4 net24
rlabel metal2 s 1610 21743 1610 21743 4 net25
rlabel metal2 s 874 21743 874 21743 4 net3
rlabel metal2 s 11914 21743 11914 21743 4 net4
rlabel metal2 s 11178 21743 11178 21743 4 net5
rlabel metal2 s 10442 21743 10442 21743 4 net6
rlabel metal2 s 9706 21743 9706 21743 4 net7
rlabel metal2 s 8970 21743 8970 21743 4 net8
rlabel metal2 s 8418 21811 8418 21811 4 net9
rlabel metal4 s 29532 22001 29532 22001 4 ui_in[0]
rlabel metal4 s 28766 22104 28826 22304 4 ui_in[1]
port 7 nsew
rlabel metal2 s 25714 20281 25714 20281 4 uo_out[0]
flabel metal4 s 31488 496 31808 21808 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 23714 496 24034 21808 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 15940 496 16260 21808 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 8166 496 8486 21808 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 27601 496 27921 21808 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal4 s 19827 496 20147 21808 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal4 s 12053 496 12373 21808 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal4 s 4279 496 4599 21808 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal4 s 30974 22104 31034 22304 0 FreeSans 600 90 0 0 clk
port 3 nsew
flabel metal4 s 31710 22104 31770 22304 0 FreeSans 600 90 0 0 ena
port 4 nsew
flabel metal4 s 30238 22104 30298 22304 0 FreeSans 600 90 0 0 rst_n
port 5 nsew
flabel metal4 s 29502 22104 29562 22304 0 FreeSans 600 90 0 0 ui_in[0]
port 6 nsew
flabel metal4 s 28796 22204 28796 22204 0 FreeSans 600 90 0 0 ui_in[1]
flabel metal4 s 28030 22104 28090 22304 0 FreeSans 600 90 0 0 ui_in[2]
port 8 nsew
flabel metal4 s 27294 22104 27354 22304 0 FreeSans 600 90 0 0 ui_in[3]
port 9 nsew
flabel metal4 s 26558 22104 26618 22304 0 FreeSans 600 90 0 0 ui_in[4]
port 10 nsew
flabel metal4 s 25822 22104 25882 22304 0 FreeSans 600 90 0 0 ui_in[5]
port 11 nsew
flabel metal4 s 25086 22104 25146 22304 0 FreeSans 600 90 0 0 ui_in[6]
port 12 nsew
flabel metal4 s 24350 22104 24410 22304 0 FreeSans 600 90 0 0 ui_in[7]
port 13 nsew
flabel metal4 s 23614 22104 23674 22304 0 FreeSans 600 90 0 0 uio_in[0]
port 14 nsew
flabel metal4 s 22878 22104 22938 22304 0 FreeSans 600 90 0 0 uio_in[1]
port 15 nsew
flabel metal4 s 22142 22104 22202 22304 0 FreeSans 600 90 0 0 uio_in[2]
port 16 nsew
flabel metal4 s 21406 22104 21466 22304 0 FreeSans 600 90 0 0 uio_in[3]
port 17 nsew
flabel metal4 s 20670 22104 20730 22304 0 FreeSans 600 90 0 0 uio_in[4]
port 18 nsew
flabel metal4 s 19934 22104 19994 22304 0 FreeSans 600 90 0 0 uio_in[5]
port 19 nsew
flabel metal4 s 19198 22104 19258 22304 0 FreeSans 600 90 0 0 uio_in[6]
port 20 nsew
flabel metal4 s 18462 22104 18522 22304 0 FreeSans 600 90 0 0 uio_in[7]
port 21 nsew
flabel metal4 s 5950 22104 6010 22304 0 FreeSans 600 90 0 0 uio_oe[0]
port 22 nsew
flabel metal4 s 5214 22104 5274 22304 0 FreeSans 600 90 0 0 uio_oe[1]
port 23 nsew
flabel metal4 s 4478 22104 4538 22304 0 FreeSans 600 90 0 0 uio_oe[2]
port 24 nsew
flabel metal4 s 3742 22104 3802 22304 0 FreeSans 600 90 0 0 uio_oe[3]
port 25 nsew
flabel metal4 s 3006 22104 3066 22304 0 FreeSans 600 90 0 0 uio_oe[4]
port 26 nsew
flabel metal4 s 2270 22104 2330 22304 0 FreeSans 600 90 0 0 uio_oe[5]
port 27 nsew
flabel metal4 s 1534 22104 1594 22304 0 FreeSans 600 90 0 0 uio_oe[6]
port 28 nsew
flabel metal4 s 798 22104 858 22304 0 FreeSans 600 90 0 0 uio_oe[7]
port 29 nsew
flabel metal4 s 11838 22104 11898 22304 0 FreeSans 600 90 0 0 uio_out[0]
port 30 nsew
flabel metal4 s 11102 22104 11162 22304 0 FreeSans 600 90 0 0 uio_out[1]
port 31 nsew
flabel metal4 s 10366 22104 10426 22304 0 FreeSans 600 90 0 0 uio_out[2]
port 32 nsew
flabel metal4 s 9630 22104 9690 22304 0 FreeSans 600 90 0 0 uio_out[3]
port 33 nsew
flabel metal4 s 8894 22104 8954 22304 0 FreeSans 600 90 0 0 uio_out[4]
port 34 nsew
flabel metal4 s 8158 22104 8218 22304 0 FreeSans 600 90 0 0 uio_out[5]
port 35 nsew
flabel metal4 s 7422 22104 7482 22304 0 FreeSans 600 90 0 0 uio_out[6]
port 36 nsew
flabel metal4 s 6686 22104 6746 22304 0 FreeSans 600 90 0 0 uio_out[7]
port 37 nsew
flabel metal4 s 17726 22104 17786 22304 0 FreeSans 600 90 0 0 uo_out[0]
port 38 nsew
flabel metal4 s 16990 22104 17050 22304 0 FreeSans 600 90 0 0 uo_out[1]
port 39 nsew
flabel metal4 s 16254 22104 16314 22304 0 FreeSans 600 90 0 0 uo_out[2]
port 40 nsew
flabel metal4 s 15518 22104 15578 22304 0 FreeSans 600 90 0 0 uo_out[3]
port 41 nsew
flabel metal4 s 14782 22104 14842 22304 0 FreeSans 600 90 0 0 uo_out[4]
port 42 nsew
flabel metal4 s 14046 22104 14106 22304 0 FreeSans 600 90 0 0 uo_out[5]
port 43 nsew
flabel metal4 s 13310 22104 13370 22304 0 FreeSans 600 90 0 0 uo_out[6]
port 44 nsew
flabel metal4 s 12574 22104 12634 22304 0 FreeSans 600 90 0 0 uo_out[7]
port 45 nsew
<< properties >>
string FIXED_BBOX 0 0 32200 22304
<< end >>
