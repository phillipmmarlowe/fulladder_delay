* NGSPICE file created from tt_um_example.ext - technology: sky130A

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VPWR VPB VNB
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

.subckt tt_um_example VGND VPWR clk ena rst_n ui_in[0] ui_in[1] ui_in[2] ui_in[3]
+ ui_in[4] ui_in[5] ui_in[6] ui_in[7] uio_in[0] uio_in[1] uio_in[2] uio_in[3] uio_in[4]
+ uio_in[5] uio_in[6] uio_in[7] uio_oe[0] uio_oe[4] uio_oe[5] uio_oe[6] uio_oe[7]
+ uio_out[0] uio_out[1] uio_out[2] uio_out[3] uio_out[4] uio_out[5] uio_out[6] uio_out[7]
+ uo_out[0] uo_out[1] uo_out[2] uo_out[3] uo_out[4] uo_out[5] uo_out[6] uo_out[7]
+ uio_oe[3] uio_oe[2] uio_oe[1]
XFILLER_0_27_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_14_161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_6_118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_8_Left_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_34_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_17_181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_37_Left_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_37_287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_12_Right_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_21_Right_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_30_Right_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_24_Left_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_27_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_6_Right_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_11_Left_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_38_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_37_288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_25_225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_0_80 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_23_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_37_289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_0_81 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_30_251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_5_111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_82 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_28_Left_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_19_Right_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_28_Right_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_37_Right_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_15_Left_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_5_112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_0_Left_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_11_147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_83 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_3_Left_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_32_Left_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_5_113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_36_281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_84 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_1_Right_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_5_114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_85 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_38_300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_15_Right_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_24_Right_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_33_Right_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_19_Left_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_5_115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_36_283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_24_220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_86 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_38_301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_21_201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_7_Left_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_22_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_36_284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_36_Left_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_20_Left_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_0_87 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_38_302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_23_Left_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_5_Right_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_36_285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_88 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_11_Right_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_20_Right_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_36_286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_33_267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_78 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_23_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_10_143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_33_268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_79 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput1 ui_in[0] VGND VGND VPWR VPWR net1 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_14_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_27_Left_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_19_190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_16_171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_9_Right_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_14_Left_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_90 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput2 ui_in[1] VGND VGND VPWR VPWR net2 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_36_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_2_Left_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_02_ _00_ VGND VGND VPWR VPWR uo_out[0] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_7_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_16_172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_8_129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_4_110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_31_Left_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_24_215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xtt_um_example_20 VGND VGND VPWR VPWR tt_um_example_20/HI uio_oe[1] sky130_fd_sc_hd__conb_1
XFILLER_0_32_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_91 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_18_Right_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_27_Right_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_36_Right_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_01_ net2 net1 VGND VGND VPWR VPWR _00_ sky130_fd_sc_hd__and2_1
XFILLER_0_20_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_19_192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_0_Right_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_27_235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_32_260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xtt_um_example_10 VGND VGND VPWR VPWR tt_um_example_10/HI uio_out[6] sky130_fd_sc_hd__conb_1
Xtt_um_example_21 VGND VGND VPWR VPWR tt_um_example_21/HI uio_oe[2] sky130_fd_sc_hd__conb_1
XFILLER_0_1_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_92 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_13_155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_182 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_18_Left_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_32_261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xtt_um_example_11 VGND VGND VPWR VPWR tt_um_example_11/HI uio_out[7] sky130_fd_sc_hd__conb_1
Xtt_um_example_22 VGND VGND VPWR VPWR tt_um_example_22/HI uio_oe[3] sky130_fd_sc_hd__conb_1
XFILLER_0_32_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_1_93 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_6_Left_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_16_175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_32_262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_35_Left_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xtt_um_example_12 VGND VGND VPWR VPWR tt_um_example_12/HI uo_out[1] sky130_fd_sc_hd__conb_1
Xtt_um_example_23 VGND VGND VPWR VPWR tt_um_example_23/HI uio_oe[4] sky130_fd_sc_hd__conb_1
XFILLER_0_20_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_14_Right_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_23_Right_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_32_Right_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_22_Left_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_16_176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_7_122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_4_Right_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_24_219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xtt_um_example_13 VGND VGND VPWR VPWR tt_um_example_13/HI uo_out[2] sky130_fd_sc_hd__conb_1
Xtt_um_example_24 VGND VGND VPWR VPWR tt_um_example_24/HI uio_oe[5] sky130_fd_sc_hd__conb_1
XFILLER_0_11_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_7_123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_32_264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xtt_um_example_14 VGND VGND VPWR VPWR tt_um_example_14/HI uo_out[3] sky130_fd_sc_hd__conb_1
Xtt_um_example_25 VGND VGND VPWR VPWR tt_um_example_25/HI uio_oe[6] sky130_fd_sc_hd__conb_1
XFILLER_0_20_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_7_124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_38_292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_4_105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xtt_um_example_15 VGND VGND VPWR VPWR tt_um_example_15/HI uo_out[4] sky130_fd_sc_hd__conb_1
XFILLER_0_11_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_10_Right_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_26_Left_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_10_Left_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_7_125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_38_293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_4_106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_26_230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_8_Right_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_13_Left_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_23_211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xtt_um_example_16 VGND VGND VPWR VPWR tt_um_example_16/HI uo_out[5] sky130_fd_sc_hd__conb_1
XFILLER_0_11_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_1_Left_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_7_126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_26_231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_23_212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xtt_um_example_17 VGND VGND VPWR VPWR tt_um_example_17/HI uo_out[6] sky130_fd_sc_hd__conb_1
XFILLER_0_31_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_19_189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_38_295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_35_276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xtt_um_example_18 VGND VGND VPWR VPWR tt_um_example_18/HI uo_out[7] sky130_fd_sc_hd__conb_1
XFILLER_0_0_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_1_89 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xtt_um_example_3 VGND VGND VPWR VPWR tt_um_example_3/HI uio_oe[7] sky130_fd_sc_hd__conb_1
XFILLER_0_37_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_38_296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_12_152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_35_277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_30_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_17_Right_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_26_Right_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_35_Right_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_17_Left_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xtt_um_example_19 VGND VGND VPWR VPWR tt_um_example_19/HI uio_oe[0] sky130_fd_sc_hd__conb_1
XFILLER_0_0_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xtt_um_example_4 VGND VGND VPWR VPWR tt_um_example_4/HI uio_out[0] sky130_fd_sc_hd__conb_1
XFILLER_0_10_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_2_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_38_297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_5_Left_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_35_278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_32_259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_32_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_34_Left_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xtt_um_example_5 VGND VGND VPWR VPWR tt_um_example_5/HI uio_out[1] sky130_fd_sc_hd__conb_1
XFILLER_0_10_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_21_Left_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_38_318 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_38_298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_3_100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_34_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_3_Right_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xtt_um_example_6 VGND VGND VPWR VPWR tt_um_example_6/HI uio_out[2] sky130_fd_sc_hd__conb_1
XFILLER_0_37_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_18_182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_38_299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_3_101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_13_Right_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_22_Right_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_31_Right_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xtt_um_example_7 VGND VGND VPWR VPWR tt_um_example_7/HI uio_out[3] sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_18_183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_6_121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_3_102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_9_Left_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_26_226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_38_Left_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xtt_um_example_8 VGND VGND VPWR VPWR tt_um_example_8/HI uio_out[4] sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_18_184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_29_246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_25_Left_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_3_103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_26_227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_7_Right_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_12_Left_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_290 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xtt_um_example_9 VGND VGND VPWR VPWR tt_um_example_9/HI uio_out[5] sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_2_94 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_29_247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_3_104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_2_95 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_18_186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_29_Right_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_38_Right_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_26_229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_31_254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_2_96 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_34_274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_29_Left_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_31_255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_16_Left_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_2_97 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_34_275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_4_Left_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_31_256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_30_Left_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_33_Left_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_2_98 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_9_135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_6_116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_16_Right_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_28_240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_25_Right_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_34_Right_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_31_257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_2_Right_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_2_99 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_20_196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_31_258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
.ends

