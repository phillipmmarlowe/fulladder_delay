magic
tech sky130A
magscale 1 2
timestamp 1709879585
<< nwell >>
rect 514 21477 31686 21798
rect 514 20389 31686 20955
rect 514 19301 31686 19867
rect 514 18213 31686 18779
rect 514 17125 31686 17691
rect 514 16037 31686 16603
rect 514 14949 31686 15515
rect 514 13861 31686 14427
rect 514 12773 31686 13339
rect 514 11685 31686 12251
rect 514 10597 31686 11163
rect 514 9509 31686 10075
rect 514 8421 31686 8987
rect 514 7333 31686 7899
rect 514 6245 31686 6811
rect 514 5157 31686 5723
rect 514 4069 31686 4635
rect 514 2981 31686 3547
rect 514 1893 31686 2459
rect 514 805 31686 1371
<< obsli1 >>
rect 552 527 31648 21777
<< obsm1 >>
rect 552 496 31808 21956
<< obsm2 >>
rect 846 507 31802 22273
<< obsm3 >>
rect 790 511 31806 22269
<< metal4 >>
rect 798 22104 858 22304
rect 1534 22104 1594 22304
rect 2270 22104 2330 22304
rect 3006 22104 3066 22304
rect 3742 22104 3802 22304
rect 4478 22104 4538 22304
rect 5214 22104 5274 22304
rect 5950 22104 6010 22304
rect 6686 22104 6746 22304
rect 7422 22104 7482 22304
rect 8158 22104 8218 22304
rect 8894 22104 8954 22304
rect 9630 22104 9690 22304
rect 10366 22104 10426 22304
rect 11102 22104 11162 22304
rect 11838 22104 11898 22304
rect 12574 22104 12634 22304
rect 13310 22104 13370 22304
rect 14046 22104 14106 22304
rect 14782 22104 14842 22304
rect 15518 22104 15578 22304
rect 16254 22104 16314 22304
rect 16990 22104 17050 22304
rect 17726 22104 17786 22304
rect 18462 22104 18522 22304
rect 19198 22104 19258 22304
rect 19934 22104 19994 22304
rect 20670 22104 20730 22304
rect 21406 22104 21466 22304
rect 22142 22104 22202 22304
rect 22878 22104 22938 22304
rect 23614 22104 23674 22304
rect 24350 22104 24410 22304
rect 25086 22104 25146 22304
rect 25822 22104 25882 22304
rect 26558 22104 26618 22304
rect 27294 22104 27354 22304
rect 28030 22104 28090 22304
rect 28766 22104 28826 22304
rect 29502 22104 29562 22304
rect 30238 22104 30298 22304
rect 30974 22104 31034 22304
rect 31710 22104 31770 22304
rect 4279 496 4599 21808
rect 8166 496 8486 21808
rect 12053 496 12373 21808
rect 15940 496 16260 21808
rect 19827 496 20147 21808
rect 23714 496 24034 21808
rect 27601 496 27921 21808
rect 31488 496 31808 21808
<< obsm4 >>
rect 938 22024 1454 22269
rect 1674 22024 2190 22269
rect 2410 22024 2926 22269
rect 3146 22024 3662 22269
rect 3882 22024 4398 22269
rect 4618 22024 5134 22269
rect 5354 22024 5870 22269
rect 6090 22024 6606 22269
rect 6826 22024 7342 22269
rect 7562 22024 8078 22269
rect 8298 22024 8814 22269
rect 9034 22024 9550 22269
rect 9770 22024 10286 22269
rect 10506 22024 11022 22269
rect 11242 22024 11758 22269
rect 11978 22024 12494 22269
rect 12714 22024 13230 22269
rect 13450 22024 13966 22269
rect 14186 22024 14702 22269
rect 14922 22024 15438 22269
rect 15658 22024 16174 22269
rect 16394 22024 16910 22269
rect 17130 22024 17646 22269
rect 17866 22024 18382 22269
rect 18602 22024 19118 22269
rect 19338 22024 19854 22269
rect 20074 22024 20590 22269
rect 20810 22024 21326 22269
rect 21546 22024 22062 22269
rect 22282 22024 22798 22269
rect 23018 22024 23534 22269
rect 23754 22024 24270 22269
rect 24490 22024 25006 22269
rect 25226 22024 25742 22269
rect 25962 22024 26478 22269
rect 26698 22024 27214 22269
rect 27434 22024 27950 22269
rect 28170 22024 28686 22269
rect 28906 22024 29422 22269
rect 795 21888 29565 22024
rect 795 19211 4199 21888
rect 4679 19211 8086 21888
rect 8566 19211 11973 21888
rect 12453 19211 15860 21888
rect 16340 19211 19747 21888
rect 20227 19211 23634 21888
rect 24114 19211 27521 21888
rect 28001 19211 29565 21888
<< labels >>
rlabel metal4 s 8166 496 8486 21808 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 15940 496 16260 21808 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 23714 496 24034 21808 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 31488 496 31808 21808 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 4279 496 4599 21808 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 12053 496 12373 21808 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 19827 496 20147 21808 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 27601 496 27921 21808 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 30974 22104 31034 22304 6 clk
port 3 nsew signal input
rlabel metal4 s 31710 22104 31770 22304 6 ena
port 4 nsew signal input
rlabel metal4 s 30238 22104 30298 22304 6 rst_n
port 5 nsew signal input
rlabel metal4 s 29502 22104 29562 22304 6 ui_in[0]
port 6 nsew signal input
rlabel metal4 s 28766 22104 28826 22304 6 ui_in[1]
port 7 nsew signal input
rlabel metal4 s 28030 22104 28090 22304 6 ui_in[2]
port 8 nsew signal input
rlabel metal4 s 27294 22104 27354 22304 6 ui_in[3]
port 9 nsew signal input
rlabel metal4 s 26558 22104 26618 22304 6 ui_in[4]
port 10 nsew signal input
rlabel metal4 s 25822 22104 25882 22304 6 ui_in[5]
port 11 nsew signal input
rlabel metal4 s 25086 22104 25146 22304 6 ui_in[6]
port 12 nsew signal input
rlabel metal4 s 24350 22104 24410 22304 6 ui_in[7]
port 13 nsew signal input
rlabel metal4 s 23614 22104 23674 22304 6 uio_in[0]
port 14 nsew signal input
rlabel metal4 s 22878 22104 22938 22304 6 uio_in[1]
port 15 nsew signal input
rlabel metal4 s 22142 22104 22202 22304 6 uio_in[2]
port 16 nsew signal input
rlabel metal4 s 21406 22104 21466 22304 6 uio_in[3]
port 17 nsew signal input
rlabel metal4 s 20670 22104 20730 22304 6 uio_in[4]
port 18 nsew signal input
rlabel metal4 s 19934 22104 19994 22304 6 uio_in[5]
port 19 nsew signal input
rlabel metal4 s 19198 22104 19258 22304 6 uio_in[6]
port 20 nsew signal input
rlabel metal4 s 18462 22104 18522 22304 6 uio_in[7]
port 21 nsew signal input
rlabel metal4 s 5950 22104 6010 22304 6 uio_oe[0]
port 22 nsew signal output
rlabel metal4 s 5214 22104 5274 22304 6 uio_oe[1]
port 23 nsew signal output
rlabel metal4 s 4478 22104 4538 22304 6 uio_oe[2]
port 24 nsew signal output
rlabel metal4 s 3742 22104 3802 22304 6 uio_oe[3]
port 25 nsew signal output
rlabel metal4 s 3006 22104 3066 22304 6 uio_oe[4]
port 26 nsew signal output
rlabel metal4 s 2270 22104 2330 22304 6 uio_oe[5]
port 27 nsew signal output
rlabel metal4 s 1534 22104 1594 22304 6 uio_oe[6]
port 28 nsew signal output
rlabel metal4 s 798 22104 858 22304 6 uio_oe[7]
port 29 nsew signal output
rlabel metal4 s 11838 22104 11898 22304 6 uio_out[0]
port 30 nsew signal output
rlabel metal4 s 11102 22104 11162 22304 6 uio_out[1]
port 31 nsew signal output
rlabel metal4 s 10366 22104 10426 22304 6 uio_out[2]
port 32 nsew signal output
rlabel metal4 s 9630 22104 9690 22304 6 uio_out[3]
port 33 nsew signal output
rlabel metal4 s 8894 22104 8954 22304 6 uio_out[4]
port 34 nsew signal output
rlabel metal4 s 8158 22104 8218 22304 6 uio_out[5]
port 35 nsew signal output
rlabel metal4 s 7422 22104 7482 22304 6 uio_out[6]
port 36 nsew signal output
rlabel metal4 s 6686 22104 6746 22304 6 uio_out[7]
port 37 nsew signal output
rlabel metal4 s 17726 22104 17786 22304 6 uo_out[0]
port 38 nsew signal output
rlabel metal4 s 16990 22104 17050 22304 6 uo_out[1]
port 39 nsew signal output
rlabel metal4 s 16254 22104 16314 22304 6 uo_out[2]
port 40 nsew signal output
rlabel metal4 s 15518 22104 15578 22304 6 uo_out[3]
port 41 nsew signal output
rlabel metal4 s 14782 22104 14842 22304 6 uo_out[4]
port 42 nsew signal output
rlabel metal4 s 14046 22104 14106 22304 6 uo_out[5]
port 43 nsew signal output
rlabel metal4 s 13310 22104 13370 22304 6 uo_out[6]
port 44 nsew signal output
rlabel metal4 s 12574 22104 12634 22304 6 uo_out[7]
port 45 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 32200 22304
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 374366
string GDS_FILE /work/runs/wokwi/results/signoff/tt_um_example.magic.gds
string GDS_START 34154
<< end >>

